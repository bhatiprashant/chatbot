id,username,user_title,raw, moderator, admin, staff, trust_level, topic_title, category_id
1143|TresataSupport||Steps to Recreate above error\n\n1. Go to Validate Step of a configured product on Pre-Prod Env\n2. Under Query Builder, Click on "Data Asset"\n3. Using the explore option create a query by adding a condition of Single equals false\n4. Click on Apply and Executed Query|false|true|true|4|Bug: Unable to Query Singleton Value|35
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
957|TresataSupport||![output_final|video](upload://9wkAkzQd1PuzMV10royH7On0iPb.mp4)|false|true|true|4|Output Full Walkthrough|87
955|TresataSupport||![Orchestrate_Final|video](upload://6bcTOYRkdzXhIKujWMKym7h0MJI.mp4)|false|true|true|4|Orchestrate Full Walkthrough|83
954|TresataSupport||![Enrich_Full_Video|video](upload://asTLKWyN4EAQ5iXMKsJs3EJ7Rl7.mp4)|false|true|true|4|Enrich Full Walkthrough|87
953|TresataSupport||![full_validate|video](upload://qsTWBSZMCEpaP4E5cPo8u2j3HIG.mp4)|false|true|true|4|Validate Full Walkthrough|86
952|TresataSupport||![trimmed_connect|video](upload://fKgFYFURX58QDTc1vWX6zjmylII.mp4)|false|true|true|4|Connect Full Walkthrough|85
950|TresataSupport||![Profile|video](upload://3xtilRJHr9ngxeK8kPW5xDaOMIN.mp4)|false|true|true|4|Profile Full Walkthrough|80
949|TresataSupport||![trimmed_prepare|video](upload://mQzU4wiHRmQGzoXtPgCplr2KGnd.mp4)|false|true|true|4|Prepare Full Walkthrough|82
948|TresataSupport||![Dashboard_Final|video](upload://5lg7mi3wS4ZIhoTyX304JuG25ky.mp4)|false|true|true|4|Dashboard Full Walkthrough|93
947|TresataSupport||![Source|video](upload://97l4dKToJMqNMmgirC9dQMToZGS.mp4)|false|true|true|4|Source Full Walkthrough|79
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
832|TresataSupport||## Azure Namespace Setup \n\nConnecting your data to our AKS cluster\n\n![Set_Up_Namespace_On_Azure|690x359](upload://kB0YXVl4JSXjaLZV0zaLEw4v08h.png)\n\nScreen: 6.0\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your Azure account. \n2. You have a storage account with Hierarchical Namespace enabled with a container inside it holding all the data you want to process. \n\n**STEPS:**\n\n1. Note down the Namespace UUID from the namespace creation panel\n2. Make sure that the storage account has "Hierarchical namespace Enabled". \n3. In the "Networking" Tab of your storage account, under "Firewall", add the address range: 0.0.0.0/0 and hit save. \n4. Create Custom Role:\n    a. In the Azure Subscription, click on "Access Control (IAM)" and click on "Add" and then "Custom Role"\n    b. Directly go to the JSON Tab and Copy Paste the following code block. Click on Review + Create\n\n```\n{\n    "id": <AUTOGENERATED_CUSTOM_ROLE_RESOURCE_ID>,\n    "properties": {\n        "roleName": "synapse-custom-role",\n        "assignableScopes": [\n            "/subscriptions/<YOUR_SUBSCRIPTION_ID>"\n        ],\n        "permissions": [\n            {\n                "actions": [\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/read",\n                    "Microsoft.Resources/subscriptions/resourceGroups/write",\n                    "Microsoft.Synapse/workspaces/read",\n                    "Microsoft.Synapse/workspaces/write",\n                    "Microsoft.ManagedIdentity/userAssignedIdentities/assign/action",\n                    "Microsoft.Synapse/workspaces/operationStatuses/read",\n                    "Microsoft.Synapse/workspaces/replaceAllIpFirewallRules/action",\n                    "Microsoft.Synapse/workspaces/operationResults/read"\n                ],\n                "notActions": [],\n                "dataActions": [],\n                "notDataActions": []\n            }\n        ]\n    }\n}\n      \n```\n\n4. Create Managed Identity:\n    a. Go to Managed Identity in the Azure portal and click on Create. \n    b. Give relevant values for the resource group, region, name, and tags and click on Create. \n5. Attach federated Credentials:\n    a. Go to the newly created Managed Identity and select federated credentials\n    b. Click on Add Credentials\n    c. Select Scenario as "Kubernetes accessing Azure Resources"\n    d. Cluster Issuer URL = "https://eastus.oic.prod-aks.azure.com/5689d11b-14df-4535-9a56-0f243ac35eca/6efda958-5385-4c8f-bc41-36ff4cac9519/"\n    e. Copy the Namespace UUID noted down from the first step - \n         Namespace = "NAMESPACE_UUID"\n    f. Service Account = "default"\n    g. Subject Identifier will be auto-filled as "system:serviceaccount::<namespaceUUID>:default\n    h. Give relevant names to the credentials\n    i. Audience = "api://AzureADTokenExchange"\n    j. Click on Add\n6. Add Role Assignments:\n    a. In that same managed identity go to the "Azure Role Assignment" and select add role assignment\n    b. Scope = Storage, Resource = <STORAGE_ACCOUNT_NAME>, Role = "Storage Blob Data Owner" and hit "Save"\n    c. In that same managed identity, again go to the "Azure Role Assignment" and select Add Role Assignment\n    f. Scope = Subscription, Subscription = <YOUR_SUBSCRIPTION_NAME>, Role ="synapse-custom-role" (This is the custom role you \n       created above. \n7. Copy the ClientID and Resource ID of the managed identity, TenantID, Storage Account Name, and Container Name to the Namespace Creation Page.\n8. After creating the namespace, the corresponding Synapse workspace will also be created with same Name as the NamesapceUUID.\n9. To give the permissions to access Synapse:\n   a. Go to the Synapse Workspace Created and click on Networking. Here add your ClientIp to the firewall and click on save.\n   b. Click on the Web URL to open the Synapse workspace and click on Manage --> Access Control --> Add Role Assignment --> Here add \n       your user as the "Synapse Administrator". (This will give you the access to add/delete role assignments.\n   c. Once you have access and you can see the other role assignments, Delete the Role Assignment for the Managed Identity as Synapse \n       Administrator.\n d. Now Add the same Role Assignment again i.e Synapse Administrator for the Managed Identity.|false|true|true|4|0.6 Set Up A Namespace On Azure|93
831|TresataSupport||## AWS Namespace Setup - Using Access Keys and Secret Keys\n\n![Set_Up_Namespace_On_AWS_Using_Access_key/Access_Secret_Key|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 5.0\n\nConnecting your data to our EKS cluster\n\n**PREREQUISITES:**\n\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n\n1. Create an IAM user and attach S3 Bucket access to that user\n    a. Go to the IAM service\n    b. Navigate to the "Users" and click on "Create user"\n    c. Give the appropriate User Name and click on Next\n    d. From the "Permissions options" select Attach Policies Directly \n    e. Click on "Create Policy"\n    f. Select JSON and paste the following in the "Policy Editor"\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    g. Review and Create the Policy and attach it to the user created in the above step\n    h. Navigate to the newly created user and click on the "Security Credentials" tab. \n    i. Click on "Create Access key" select "Command Line Access" and check on the confirmation button\n    j. Download and open these keys and paste appropriate values for AccessKey and SecretKey in the Create namespace page.\n\n---\n**NOTE**: Substitute these values appropriately in the JSON\n* S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to.\n\n* NAMESPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page.\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n---|false|true|true|4|0.5 Set Up A Namespace On AWS Using Access Key/ Secret Key|93
830|TresataSupport||# AWS ROLE ACCESS\n\n![Set_Up_Namespace_On_AWS_Using_Role_ARN|690x359](upload://xH69vv1YISaUPy9LlUQjo0WaISF.png)\n\nScreen: 4.0\n\nConnecting your data to our EKS cluster (Recommended method)\n\n**PREREQUISITES:**\n1. You (ADMIN) have administrator-level privileges in your AWS account. \n2. You have an S3 Bucket where the data is stored\n\n**STEPS:**\n1. Note down the Namespace UUID from the namespace creation panel\n2. In your AWS Account, create an Identity Provider:\n    a. Go to the IAM service\n    b. Navigate to the "Identity Providers" and choose "Create Provider"\n    c. Select "OpenID Connect" as the provider type.\n    d. Provider URL = "https://oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n    e. Click on Get thumbprint and AWS will generate this value. \n    f. Audience = "sts.amazonaws.com"\n    g. Review the information and then click on "Add Provider"\n3. Create an IAM role and Trust relationship so that only the Namespace created by you, will have access to data\n    a. Go to the IAM service\n    b. Navigate to the "Roles" and select "Create Role"\n    c. Select Custom Trust Policy and add this JSON\n\n```    \n{\n    "Version": "2012-10-17",\n    "Statement": [\n        {\n            "Effect": "Allow",\n            "Principal": {\n      "Federated": "arn:aws:iam::<YOUR_ACCOUNT_ID>:oidc-provider/oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550"\n            },\n            "Action": "sts:AssumeRoleWithWebIdentity",\n            "Condition": {\n                "StringEquals": {\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:sub": "system:serviceaccount:<NAMESPACE_UUID>:default",\n                    "oidc.eks.us-east-1.amazonaws.com/id/E1B2EB40F8031126E7E6AA1D69937550:aud": "sts.amazonaws.com"\n                }\n            }\n        }\n    ]\n}\n```\n   - d. To attach the policy to the role, select "Create Policy" and add this JSON:\n\n```\n{\n    "Statement": [\n        {\n            "Action": [\n                "s3:GetBucketLocation",\n                "s3:ListBucket"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<S3_BUCKET_NAME>"\n        },\n        {\n            "Action": [\n                "s3:GetObject",\n                "s3:GetObjectTagging",\n                "s3:PutObject",\n                "s3:DeleteObject",\n                "s3:ListMultipartUploadParts",\n                "s3:AbortMultipartUpload"\n            ],\n            "Effect": "Allow",\n            "Resource": "arn:aws:s3:::<s3_BUCKET_NAME>/*"\n        },\n        {\n            "Action": [\n                "athena:StartQueryExecution",\n                "athena:GetQueryExecution",\n                "athena:GetQueryResults",\n                "athena:StopQueryExecution",\n                "athena:ListQueryExecutions",\n                "athena:CreateWorkGroup",\n                "athena:GetWorkGroup"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:athena:us-east-1:<YOUR_ACCOUNT_ID>:workgroup/<NAMESPACE_UUID>"\n            ]\n        },\n        {\n            "Action": [\n                "glue:GetTables",\n                "glue:GetTable",\n                "glue:CreateTable",\n                "glue:UpdateTable"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:table/<NAMESPACE_UUID>/*"\n            ]\n        },\n        {\n            "Action": [\n                "glue:CreateDatabase",\n                "glue:GetDatabases",\n                "glue:GetDatabase"\n            ],\n            "Effect": "Allow",\n            "Resource": [\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:catalog",\n                "arn:aws:glue:us-east-1:<YOUR_ACCOUNT_ID>:database/<NAMESPACE_UUID>"\n            ]\n        }\n    ],\n    "Version": "2012-10-17"\n}\n```\n*\n    e. Give this policy an appropriate name and attach it to the role you are creating. \n    f. Give this role an appropriate name and click on "Create Role"\n    g. Copy the RoleArn of this role and paste it under the roleArn box in the "Create a Namespace" page.\n\n---\n**NOTE**: You need to substitute these values appropriately in the JSON\n\n* YOUR_ACCOUNT_ID - This is your AWS subscriptions Account ID. You will get this information if you click on your user in the upper right-hand corner of your AWS Console.\n\n* NAMESCPACE_UUID - This is the value you noted down in the very first step. Copy and paste the value from the Namespace Creation Page. \n* YOUR_S3_BUCKET_NAME - Paste the S3 bucket name of the bucket you are giving us access to. \n---|false|true|true|4|0.4 Set Up A Namespace On AWS Using Role ARN|93
806|TresataSupport||\nNow that you have successfully connected to our namespace, now its time to start the first product on TRESATA. In this post let's see how to create a new product from your dashboard, how to edit them if required and many more. So with no further ado, let's begin.\n\n**STEPS TO ADD NEW PRODUCT**\n\n![Dashboard_Create_New_Product|690x359](upload://1ZUIc2JBUcjqykts1QvWWTLFqkE.jpeg)\n*Screen:3.0*\n\n![image|690x347](upload://pbDMP5koh3fLMbfmKWQbYsU0PrY.png)\n*Screen 3.1*\n\n![Dashboard_Add_Name_Description|690x359](upload://6W3sc22HR6e09e4Zf8djFBlo1Kl.jpeg)\n*Screen: 3.2*\n\n* For admin users, they can easily get started off with creating their product simply just clicking on the *Create Product* button as shown in the screen 3.0\n* Next choose a category from the list above to select product type. You can choose NOTA(None of the above) when they want to give custom category. These categories becomes prominent as TRESATA will suggest customised cleaners and resolution logic for your product.\n* After which a pop-up comes for you to provide a name for your product and a small description about it as shown in screen 3.1. After which it takes the you to the Sourcing Step.\n* If you are not an admin, and just received link to sign up to the product, then you will have to wait for your admin to approve your namespace. Only approved users are allowed to create their products. So be sure to ping your admin if not approved yet.\n\n---\n**EDIT PRODUCT NAME**\n\n![Dashboard_Edit_Product|690x359](upload://qTkS0gJzWVg5lRFxLohRk5Y7fKy.jpeg)\n*Screen: 3.2*\n\nIn the Screen 3.2, as you can see the list of products that has been created in this particular account or you can say in the namespace. If you want to edit the name or the description of the product, you has to simply click on the *edit icon* as seen above.\n\n![Dashboard_Naming_Best_Practice|690x359](upload://1XSsuWCUOCCP54Tp0SBDFaeWrKL.jpeg)\n*Screen: 3.3*\n\nThe name of the product can not have any special symbols or product names can not be repeated in the given namespace.\n\n---\n**Go to Step in Product Listing**\n \n![Dashboard_Product_Stage_Listing|690x359](upload://4OIRI6jcrQSbFiRkHwtQVRqiW8v.jpeg)\n*Screen: 3.4.1*\n\n![Dashboard_Product_Stage_Listing_updated](upload://dfwyzahbmoOfPIcbpNvKKlUzKbN.jpeg)\n*Screen: 3.4.2*\n\nIf the product has been created, and some steps of TRESATA has been finished. In that case, you can directly access that step with the help of a drop-down to view or continue working from that step directly As seen above in Screen 3.4.1, choose any of the steps that has been listed, and clicking on the button *GO* will take us to corresponding home-screen immediately \n\n----\n\n**DELETE PRODUCT**\n\nProducts can be deleted easily from the Dashboard with the delete option that is present next to edit button. If you are an Admin, then you will get couple of extra features to handle the deleted products. \n\nMore information on Admin rights of Deleted product was discussed in the previous post  [here](https://community.tresata.com/t/2-admin-panel-actions/566). \nFeel free to check them out. Let's begin our first step of your Data transformation which we call as Sourcing in the next post.. See you soon.!!|false|true|true|4|0.3 Create a new Product|93
801|TresataSupport||As we have started off with the first step to use product TRESATA by initial sign up process and login. It is important to note that there are few privileges that is availed only to an Admin user. This post is aimed to list down them together so that your product can be managed effectively.\n\n**MANAGE NAMESPACE**\n \nNamespace plays a very important role for our product, without which we wont be able to connect to our data. Hence handling it better becomes crucial.  When an admin user subscribes product TRESATA, soon after the payment completion they will be taken to the TRESATA Admin Panel. So the screen 2.0 shows how  *Admin Panel* looks like. \n\n**Namespaces:** \n\n![Admin_Panel_Screen|690x359](upload://xcCloyhnnEkdiKo5T2DiAA0SOu3.jpeg)\n*Screen: 2.0*\n\nThis tab shows the details of your namespace. Name of the namespace that was created during the sign up process will be shown here as seen in Screen 2.0\n\n----\n\n**Products:** \n\n![Admin Panel-Add_Product|690x359](upload://mzNDtWVUhiiRGZ4pIYvvrpJQsLP.jpeg)\n*Screen: 2.1.1*\n\n![Admin Panel_Add_Product|690x358](upload://kfVDTqTcYgUcGxmYNp3EgOovUXW.jpeg)\n*Screen: 2.1.2*\n\nOnly admin user can create products from the Admin Panel screen, and assign users to it. Admin will have to click on the Products Tab to add a new product as shown in Screen 2.1.1.  Admin has to enter Product Name, with a small Description and Users to that Product. As seen in the Screen 2.1.2, Admin can simply choose their users from the drop down list.\n\n**Note**: \nOnly one user can be assigned to every product. Admin can create multiple products but each product shall have just one user handling it. \n\n**PRODUCT ACTIONS**\n* **Edit:**\n\n![Admin Panel_Edit_Product|690x359](upload://rsuG8LHePFFmbQfuRf8JB5VGhp7.jpeg)\n*Screen: 2.2*\n\nAdmin can change the Name and the Description of the product anytime according to their requirement. Once a User has been assigned to a product, that can not be changed under any circumstances. So it's important to the Admin to be cautious while assigning Users to their product. \n\nThere will be an upgrade very shortly allowing users to  collaborate with their co-data engineers, so stay tuned..!!!\n\n* **Delete:**\n\n![Admin Panel_Delete_Product|690x359](upload://qtIhNy62C5dwIr1ZF1f1csU9y4f.jpeg)\n*Screen: 2.3*\n\nAdmin can also delete their products easily by clicking on the delete button as shown in the Screen 2.3\n\n![Admin Panel_Select_Multiple_product|690x359](upload://osyveTf1jMPI16wASQ3hMSDFtR2.png)\n*Screen: 2.4.1*\n\n![Admin Panel_Delete _All|690x359](upload://baoqkaJfDxnFsBl5CTNWRGnlHWn.png)\n*Screen: 2.4.2*\n\nAdmin can also delete multiple products together by selecting them with the checkbox shown in the Screen 2.4.1 and then continuing to delete all as seen in 2.4.2\n\n----\n**Users:** \n\n![Admin Panel_Add_Users|690x359](upload://7WBpzAmQhxg84581LrV3dIGGWir.png)\n*Screen: 2.5*\n\nOnly Admin user will be able to add new users to the namespace that they just created. In order to do so, click on the tab of Users, hit on the button *Add Users* as seen in Screen 2.5\n\n![Admin Panel_Add_Recipients_email|690x359](upload://kACKMdJp88uhqxp6nulmThhPLcu.jpeg)\n*Screen:2.6*\n\nAdmin then has to add the email of the list of user they wish to add in the namespace\n\n![Admin Panel_Users_List|690x359](upload://byZ2E8lXs6ns2s03uzauXnLfzGs.jpeg)\n*Screen: 2.7.1*\n\n![Admin Panel_Invites_Sent|690x359](upload://q2EQrSYkfAQzMtOvBlnrUVi6dZt.png)\n*Screen: 2.7.2*\n\nAs shown in the Screen 2.7.1, even multiple users can be added by Admin to send invites to join the product. Soon after clicking on the button Send Invites, a email will be sent to every user to join TRESATA.\n\n**IMPORTANT NOTE**\n\n1. When user accepts the invite, the status of the User turns from red tag *Pending* to  green tag *Accepted*\n2. When users join through the invite sent by Admin, after user login, next Admin has to also approve them to join the Namespace too. If not, then users can not create any products on TRESATA\n\n----\n\n**CONSUMPTION**\n\n\n![image|690x325](upload://orjOxekPrmDxvRCkFEatLIDkdhE.png)\n\n*Screen: 2.8*\n\nAdmins can keep track of the CPU consumption and  Billing cost for the selected period of time as seen in above. User can also view details of avg and max consumption of CPU units and Billing cost when they hover over the graph.\n\n----\n**DELETED PRODUCTS**\n\n![Admin Panel_Deleted_Products_list|690x359](upload://wESaTWb2yTFHKIXSvnmwqNTi5vB.jpeg)\n*Screen: 2.9*\n\nThis feature is available only to an Admin User. So under the Tab of Deleted Products, users can find a list of all products that was deleted by them and deleted by the users that they assigned.\n\n![Admin Panel_Restore_Option|690x359](upload://85JfHdtCNQkWQMt2jAKUkoAYgRM.jpeg)\n*Screen: 2.10.1*\n\n![Admin Panel_Delete_Forever_Option|690x359](upload://idZjx9E0QTbVYB2DC8dWcbejWz.png)\n*Screen: 2.10.2*\n\nThe users can either restore the deleted product, which will again reflect back in the deleted users environment, or to delete it permanently, click on the button called *Delete Forever* to get them out of your namespace completely.\n\n![Admin Panel_Mass_Action|690x359](upload://6iYKh27n1pTRf4jneEAX1Q8s0qN.png)\n*Screen: 2.11*\n\nThe above screen the representation of how we can restore or delete multiple deleted products.\n\nThis is the overall walk through on Admin Panel, more details to get started with your first product is coming soon in the next post. \n\nSo stay Tuned...!!|false|true|true|4|0.2 Admin Panel Actions|93
800|TresataSupport||**Introduction**\n\nWelcome..!! Excited, as we take the first step towards an incredible journey of discovery, transformation and enrichment. This is the place for you all to unlock the power of data to enrich life.\n\nBut before we dive in, let's start with the first step which is signing up to our product **TRESATA**. This post is aimed to help you to get started with the seamless sign up process.\n\n**Steps To Sign Up:**\n\nYOU will be able to join TRESATA product from the Tresata website, with the three options to get started, which are :\n**Try for Free**, **Upload** and **Access**\n\n![image|690x349](upload://uXD7N0toDUZdkBXdc8swg6NdSZ8.png)\n *Screen: 1.0*\n\nClick on **Try For Free**, if you want to use our product and playaround using pre uploaded tresata files. \nClick on **Upload**, if you want to upload your files in Tresata's storage account and get started with the product.\nClick on **Access**, where you can link your cloud storage with the Tresata.\n\n**Environment Selection:**\n\n![image|690x346](upload://1LFAQYo45TqcColku3E6j5ch7uY.jpeg)\n*Screen: 1.1*\n\nYou are given with two options as you can see on the Screen 1.1. According to the requirement of the environment, you can choose either AWS or Azure. The sign up process vary a little based on the kind of choice is made\n\n**User Information:**\n\nThe next step is to complete sign up process by providing essential information:\n\n\n![Sign_Up|690x391](upload://r7vDq8kCO6kCeehRb4Cn67iEpFL.jpeg)\n*Screen: 1.2*\n\n* Name\n* Email\n* Password (with specific criteria)\n* Confirm Password\n* Checkbox to agree to our terms and conditions.\n* You can review our terms of service by clicking on the provided link.\n\n**Verification Email:**\n\n![image|676x500](upload://g4eE8Mubn5AkEfhWwEzidb1M869.png)\n\n*Screen: 1.3*\n\nOnce you hit the sign-up button, you will receive an email with a verification code along with a login link. This is for two-factor authentication to confirm your account.\n\n**Setting Up Your Namespace:**\n\nAfter confirming your account, you'll need to set up a "namespace." The process differs depending on your chosen environment:\n\n**AWS**: \n\n![AWS_Namespace|690x359](upload://aT29DpSvk5M9tehF0WThujPxgqZ.png)\n*Screen: 1.4*\n\nYou'll be prompted to provide:\n\n* Namespace alias name: Need to be unique and also an error message will guide you if it already exists\n\n* Role ARN: If you choose to set up your AWS account using a Role ARN (Amazon Resource Name), you need to provide the Amazon Resource Name of the IAM role that TRESATA will assume. This role should have sufficient permissions to access the necessary AWS resources.\n\n* Access Key and Secret Key: If you opt for the Access Key and Secret Key method, you'll need to provide:\n\n* Access Key: This is a unique identifier used to authenticate with AWS services.\n* Secret Key: This key is used as part of the authentication process along with the access key.\n\n* Configure AWS S3 Bucket: You need to specify the details of the AWS S3 bucket where your data sources are stored. This typically involves providing the:\n\n* Bucket Name: The name of the AWS S3 bucket.\n\n* For all the first time users, we have a detailed document on steps to create your namespace on AWS   [click here](https://docs.google.com/document/d/1zR67Hjo2jbH_kii2kZc-C5m8sq12T0ogn_5nt4P0HF4/edit)\n\n**Azure**: \n\n![Azure_Namespace_Setup|690x359](upload://fi1HNPBKI4LGoSKhUVDsbTMfWSd.png)\n*Screen: 1.5*\n\nYou'll be prompted to provide:\n\n* Namespace Alias Name: Provide a unique name that will serve as an alias for your namespace. This is what you'll use to reference your namespace within TRESATA. If the name is already in use, you'll receive an error message and will need to choose a different name.\n\n* Namespace Key: An auto-generated alphanumeric key will be provided to uniquely identify your namespace. This key is crucial for secure access to your namespace and TRESATA resources.\n\n* Azure Account Details: To connect TRESATA with your Azure account, you'll need the following information:\n\n* Client ID: This is the unique identifier for the application or service principal in Azure Active Directory that TRESATA will use to access Azure resources.\n\n* Tenant ID: This is the identifier for your Azure Active Directory tenant.\n\n* Storage Account Name: The name of the Azure Storage Account where your data sources are stored.\n\n* Container Name: The name of the container within the Storage Account where your data resides.\n\n*  For all the first time users, we have a detailed document on steps to create your namespace on Azure, [click here](https://docs.google.com/document/d/1ytCZ33m-jErwmrU5JL4sj2C997350pjfkrphkib-7d8/edit?usp=sharing)\n\n**Logging In:**\n\n![User_Log_in|690x391](upload://4JIZac164jREDp2hLR4f2HP3mkJ.jpeg)\n*Screen: 1.6*\n\nOnce user has  successfully signed up and confirmed your account, you'll land on the welcome login page. Here's what you need to know about the login process:\n\n* Provide users registered email and password to log in.\n* If you've forgotten your password, we offer a password recovery option.\n* New users who haven't signed up can use the provided link to join the TRESATA platform.\n* Once you log in, you can start exploring and utilising the TRESATA product.\n\n**Forgot Password**\n\n![Login_Forgot_Password](upload://uybDyuyLaFecitCb98SwdxPVohd.jpeg)\n*Screen: 1.7.1*\n\n![Login_Reset_Forgot_Password](upload://nWtttmT9SOiNQp2AWKajPCJJs69.jpeg)\n*Screen: 1.7.2*\n\nForgot your password ? Never-mind, we have got you covered. Just click on the forgot password option, and provide the username as shown in the Screen 1.7.1, and then you will be getting an automated reset password link on their mail list. Simply click on it and a Screen 1.7.2 will appear to reset and confirm your new password. And so, you're all set to access TRESATA..!!!|false|true|true|4|0.1 Sign Up for TRESATA|93
796|TresataSupport||This category consists of all the relevant steps for getting you started on using our product TRESATA\n\n* https://community.tresata.com/t/0-1-sign-up-for-tresata/565?u=tresatasupport\n* https://community.tresata.com/t/0-2-admin-panel-actions/566?u=tresatasupport\n* https://community.tresata.com/t/0-3-create-a-new-product/571?u=tresatasupport\n* https://community.tresata.com/t/0-4-set-up-a-namespace-on-aws-using-role-arn/584?u=tresatasupport\n* https://community.tresata.com/t/0-5-set-up-a-namespace-on-aws-using-access-key-secret-key/585\n* https://community.tresata.com/t/0-6-set-up-a-namespace-on-azure/586?u=tresatasupport\n* https://community.tresata.com/t/dashboard-full-walkthrough/667?u=tresatasupport|false|true|true|4|About the Admin category|93
795|TresataSupport||**Getting Started with Output**\n\n![Enrich_Output_Home_Screen|690x359](upload://2tRSwTT7MfLw6b7M64EOeILmLRa.png)\n*Screen: 2.0*\n\nAs shown in Screen 2.0, from the list of Output sources, users are given two choices to select their Output data\n\n1. **Universal (Per Data Source)**:\n\n![Enrich_Universal_Output|690x359](upload://7UXxIpD3l3SEMtl5afk2adYXm0k.png)\n*Screen: 2.1*\n\nThe Screen 2.1 shows the usage of Universal Output. In this method, users are given the option to customize the output schema for every data source. \n\n* **Raw Data** is your initial sourced data\n* **Cleaned Data** is the data after we finished data cleaning in Prepare Step\n* **Enriched Data** is the data after applying optimal rules to get Golden Records\n\nWith the above 3 options, users can select the required schema simply by clicking on the checkbox next to it as seen in Screen 2.1. The schema is source dependent and different schema can be selected for every data source\n\n2. **Enriched**:\n\n![Enrich_Enriched_Output|690x359](upload://d4EQS0XzASYtJUbpiMjGm1FTcym.png)\n*Screen: 2.2*\n\nAs seen earlier in the Universal Output step, the same process is followed for Enriched Output too. The main differentiator between the two is that one output schema will be generated for all the Data Sources forming a standardized global output. And Raw Data fields can not be considered for Enriched Output. \n\nUsers can select any schema that they wish to view output for and click on the button *Initiate Output* to get your Final Output.|false|true|true|4|6.2 Final Output|87
794|TresataSupport||One of Tresata's core capabilities is Enrich, allowing you to choose the best, most accurate values to create a *golden record* for each of your TresataIDs as well as tailor the output files to best feed downstream usage.\n\nThis post will provide high level information on why Enrich is important and it will briefly discuss its capabilities.\n\n**GOLDEN RECORD**\n\nHaving assigned TresataIds (TIDs) to records, you can now filter for a TID to view all the records describing one entity. However, what if you wanted to create one record, including the best, most accurate information for all of the available fields? That can be done using the Enrich feature.\n\n**STEPS TO SELECT YOUR ENRICH FIELDS**\n\n![CLick_On_Initiate_Enrich|690x359](upload://pGK0Cwne78QDwgoNmGPi1k99Ui2.png)\n*Screen: 1.0*\n\nBefore we start to choose fields for our Golden Record, it's important to shed light on a few sets of rules upon which the best fields can be selected by the user. In the Enrich stage, there are two main categories of enrichment logic available (Table and Field Preferences) and can all be configured via drag and drop operations.\n\n\n1.**Field Preferences**:\n\n![Enrich_Select_Canonical_Field|690x359](upload://eT5VFmsUAOFRbze67Q0QWS5oy8s.png)\n*Screen: 1.1*\n\nThis category will allow you to select the best value for a field to populate your Golden Record.  To use this rule, the user has to first select a Canonical Field, on the left side bar as seen in Screen 1.1. \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.2*\n\n* **Expression:** As seen in above in the Screen 1.2, by selecting this option, users can specify custom logic for how to identify the best information for this field. Expression allows you to pick a value coming from a record that meets specific ranking criteria on a field of your interest. Notice the following example:\n\n*While gathering information for all the bookings by *\n\n\nTaking the example of *FunAirways* from before,  Prefer First name on the expression of Create Date. So the system will set Best First Name based on the latest Create Date value.\n\n![Enrich_Count_Preference|690x359](upload://8YEE2O4FHyZEvXJI0UBXOEbY3xR.png)\n*Screen: 1.3*\n\n* Count: This option allows the user to select a particular field on the basis of the most frequent value. A counting algorithm is run in the background on the selected canonical field values. Continuing from the example above, Prefer First Name on the count of Tickets booked. \n---\n2.**Table Preferences**: \n\n As the name suggests this category is used by users to choose a source as the best information for the Golden Record. We can further see 2 ways to choose best dataset.\n\n![Enrich_Prefer_Data_Set|690x359](upload://pvOxebvRcW7PVOCyODN19re1s4P.png)\n*Screen: 1.4*\n\n* **Prefer:** Selecting Prefer Rule is simply telling Tresata, that the selected data source is the most trusted source. Now our algorithm will assign high scores on the preferred sources and choos its field values for all the canonicals from that preference.  \n\n![Enrich_Rank_Records|690x359](upload://8ZqZSNBsm7pYzc0WzJp3jsGBrIh.png)\n*Screen: 1.5*\n\n*  **Rank:** Just giving a preferred data source might not be enough when users are dealing with complex data. So to facilitate that, there is another option called RANK. Here users can choose Rank as a criteria to sort their best data, so that those fields get prioritized. In the Screen 1.5, as you can see, users can select any canonical from the available list. Users can give their preferences by allocating a specific rank to it.\n\n---\n![Enriched_Profile_Heat_Map|690x359](upload://bBtvdWZ4WaClfitzHqnva5vOMXF.png)\n*Screen: 1.6*\n\nTo make sure you are applying the right logic to select your Golden Record, users can also make use of the profiled Heat map to understand data quality and get accurate canonicals for enrichment.\n\n![Enrich_Initiate|690x359](upload://l6T637D8IlyyiQBodf80uWebED0.png)\n*Screen: 1.7*\n\nWhen user finalizes their enrichment logic, it is good to initiate the enrich step to apply all the selected rules. Users will be allowed to add any number of rules that suites their use case. Users can also edit and delete rules before clicking on the button *"Initiate Enrich"*\n\nThis will now create Optimal Output values that contain Golden Records with the best attributes.\nIn the next post, let's view the final transformed data.|false|true|true|4|6.1 Enrich & Its Significance|87
789|TresataSupport||**** \n\nIn the previous post, the importance of Validate as a step was discussed, and the main terminology and features explained. However, there is more to investigating Connect results and identifying areas for improvement: it takes investigation and evaluation of findings to pinpoint what is wrong when it comes to your Connect configurations.\n\nThat's why this post will walk you through how to evaluate and understand your Validate metrics and where to look to find some of the most common resolution gaps.\n\n**OVERALL STATISTICS**\n\nAs discussed on the earlier post, one of the main metrics provided throughout the Validate steps are the overall statistics on the top of the *Data Products Statistics* panel (*screen 1.0 below*).\n\n![Screen Shot 2023-08-20 at 3.34.18 PM|690x359](upload://6AHtYe11wsAZK5hDyMhCF74Y4Pf.png)\n*Screen 1.0*\n\nAs shown above, those statistics include:\n\n* \\# of Tresata IDs (TIDs)\n* \\# of Records\n* \\# of Data Sources\n* Avg. # of Sources per TID\n* Avg. # of Records per TID\n* Singletons\n* Spanning\n* Trapped\n\nAll the above are aggregated across all your sources, giving you a quick overview of everything within your data. But how should they be evaluated?\n\nTo begin with, the overall ***# of TresataIDs*** can show you how many entities have been identified within your data (i.e. how much your records have compressed). A very low number of TIDs compared a very high number of records can indicate over compressing ("loose" restrictions on what should bring records together). On the other hand, having too many TresataIDs can be a sign of undercompression (very restrictive connect logic) where records that should have connected don't. Of course, how much compression should be expected is relative to your use case. Let's look at the two following FunAirways use cases:\n\n* *As a data scientist at FunAirways, I am looking on all of the bookings with us for flights from the Charlotte airport by our loyalty clients (the ones signed up for our loyalty program, flying frequently with FunAirways). As I am trying to identify **how many clients** have booked with us, I am not interested on the number of bookings but rather, the unique number of clients that made them. Thus, as one client makes multiple bookings throughout a year, I should expect a low number of TIDs in relation to the number of records (number of bookings).*\n\n* *As a data scientist on FunAirways marketing team, I am trying to identify how many clients have signed up on your loyalty promotional program. For that, I am looking through the loyal customers dataset, which includes the names of the loyal customers and the unique key assigned to them by us upon sign up. On such a use case, compression is expected to be low as no customer is allowed to sign up for the promotional program twice and thus, duplication is unexpected. So, I would expect a high number of TIDs, relative close to the number of records...*\n\nSimilar way of thinking should be applied to statistics like the **Avg # of Records mer TIDS**. However, statistics like **Singletons, Trapped** and **Spanning** have some more interesting insights. As explained on the last post\n\n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn’t connected with any other record.\n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source.\n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s).\n\nAs it can be derived, the closer to 1:1 the ratio is between records and TIDs, then higher the number of Singletons will be. Similarly, the more compression we are seeing, the highest the number of Trapped and Spanning will be. But, there is more to be derived from such statistics:\n\n* *As a data scientist in FunAirways, I am trying to identify how often customers book tickets but don't actually check in for their flights. For that use case, I'll use my *booking* and *ticketing* data sources. In theory, each record in booking should connect against a record in ticketing as usually, people that book a flight eventually check in for it too. In such a use case, I should expect a high number of Spanning TIDs (TIDs with records across different sources) as it would be an unusual case to have a customer who booked a ticket but didn't check in (and eventually missed the flight).* \n\n**DATA INTEGRITY CHECK**\n\nAll the above findings, while applicable on an overview level, they are also important when looking at each source separately as, with a more granular view, you are able to pinpoint the error more accurately.\n\nNow, rather than looking at those across sources, the user can identify if there is over compression or under compression within a source, which can help when investigating what part of your Connect logic has caused the incorrect resolution. Imagine a scenario where one source has unexpected high average records per TID. While that can be tricky to identify if you have many more sources on your Data Product, especially as they interact with each other, it becomes much clearer when separating those statistics on a source level.\n\n**CROSS-DATA SOURCE OVERLAPS**\n\nAnother interesting metric, besides how many records have connected, is how many of those have connected across what data sources. As showcased above, there is different expectation on how much records should connect within or across sources, based on the information they have. Knowing what's expected it (based on your business logic) can be very valuable when evaluating overlap statistics. \n\nSource overlaps are very useful to show how your records have connected, what sources have the highest overlaps and more. Notice on screen 1.1:\n\n![Screen Shot 2023-08-20 at 4.31.41 PM|690x359](upload://xztvJCYMHw8RjV93RhpDsmNCdV3.png)\n*Screen 1.1*\n\nOn the table s on the screen, you can find the exact resolutions metrics for each data source permutation set that records have connected. Based on the table, 56% of all the records belong to a TID that only spans two sources, ***finance*** and ***esg***. Based on your domain knowledge, those statistics can either validate what you initially expected or point you to the source of the problem.|false|true|true|4|5.2 How To Validate Your Results|86
788|TresataSupport||At this point, records from each siloed source are connected with each other, using a tresataId to identify entities rather than records. Having connected your data, the next step is to investigate the accuracy of your resolution and identify areas of improvement. This post will:\n\n* Explain what is the Validate step and why it is important for an accurate Data Product\n* List and briefly describe its most important features\n\nLet's dive right in...\n\n**WHAT IS VALIDATE**\n\nValidate is the next step right after configuring Connect. In terms of user actions, Validate is automatically kicked off after successful completion of the Connect job, and upon completion if provides you with important metrics to evaluate the performance of your Connect logic. All in all, it is a hub of statistics and metrics, available in tabular format as well as a *csv* export report. \n\nAll the above are interesting, but...\n\n**WHY IS VALIDATE IMPORTANT**\n\nAccurate resolution is an outcome of an iterative process, where you configure, validate the output and adjust your logic until you get optimal results. On that cycle, Validate holds a crucial role as it provides visibility on how good your Connect output is. Without the Validate statistics, identifying resolution gaps and tuning your logic would be impossible and thus, accurate Data Products would be much more difficult to achieve. \n\n **MOST IMPORTANT FEATURES**\n\nTresata's Validate statistics suite comprises of various level of metrics, from overview statistics all the way to source specific ones. However, before focusing on what those are, it's important to understand some key terminology that will be referenced in the Validate section:\n\n* **Overcompression**: is the concept of forcing too many records to link with each other, often causing incorrect connections, bringing together records that should be separate. It is often caused by "loose" Connect logic, where the user isn't strict enough on what should link two records together. \n* **Undercompression**: is the concept of missing out on connections between records. It leads to incomplete or fragmented data connections, leaving records separated when they should have connected. This can result in lost insights and a less comprehensive view of the data landscape and it can be caused by very restrictive Connect logic. \n* **TresataID**: a unique identifier used to identify entities across many records & sources. In other words, when records connect with each other during Connect, they will receive the same tresataId, which then can be used to identify all the records related to the same entity. \n* **Singletons**: are tresataIds assigned to one record only. In other words, that record hasn't connected with any other record. \n* **Trapped**: are tresataIds that connect records from one source only. In other words, the records with that tresataId have connected only with records within the same source. \n* **Spanning**: are tresataIds that connect records across many different sources. In other words, the records from that tresataId have connected with records from different source(s). \n\nHaving explained those important concepts, let now take a quick look on Validate's metrics that will enable you on your investigations:\n\n* **Overview stats**: will include statistics such as *# of tresataIds*, *# of Records*, *# of Data Sources*, *Avg. # of Sources per TID*, *Avg. # of Records per TID*, *Singletons*, *Spanning*, *Trapped*. \n* **Counts per Data Source**: will include most of the metrics above for each data source, to provide an extra layer of granualarity.\n* **Cross-Data Source Overlaps**: will include *Data Source Combinations*, *# of Records* and *% of Records Overlapped*. This metric will show how many records overlapped (connected) between sources and what is that percentage compared to all of the connections. \n\nThe above metrics are a starter pack on identifying areas of improvements on your connection logic. Checkout the next post for a deep dive on how to utilize them to improve the efficiency of your Connect step!|false|true|true|4|5.1 Validate & Its Significance|86
780|TresataSupport||**SUMMARY**\n\nRegular Expressions or RegEx, are a powerful feature when it comes to cleaning data, aiding in the filtration and substitution of different data patterns. In addition to all the cleaners that Tresata offers, this post will help users fully harness the capabilities of Regex-Filter functionality\n\n\n**LIST OF COMMONLY USED REGEX FILTER  EXPRESSIONS**\n|Name|Regex Expression|Description|Example|Output\n|---|---|---|--|--\n|Accept Numbers | ^[0-9\\]+|Accepts only characters from 0 to 9 and '+' sign indicates to accepts all digits entered|12345|12345\n||||ab123| None\nExclude Special Characters|^[A-Za-z0-9\\]+$|Matches with characters A to Z, a to z and 0-9|hello123| hello123\n||||hello@me| None\nAccept Valid Email ID|^[a-zA-Z0-9._%+-\\]+@[a-zA-Z0-9.-]+\\\\.[a-zA-Z]{2,}$| [A-Za-z0-9\\_] represents characters from a to z with 0 to 9 digits. '@' sign is a must to validate the regex followed by any characters from a to z in lowercase then comes '.' a period with a to z characters again|user@gmail.com | user@gmail.com\n||||user@gamil|None\nPhone Number Validator|^[+\\]{1}(?:[0-9\\\\-\\\\(\\\\)\\\\/\\\\.]\\\\s?){6,15}[0-9]{1}$|Accepts any country code with the condition of starting with a plus sign (+) and then checks for 10 digits in the phone number|+1 7878 123456 | +1 7878 123456\n||||+1 7875 1234 | None\nCredit Card Validation|^(\\\\d{13,16})$|Accepts 13-16 digits of numbers shows none, if this condition is not satisfied| 1234567890123345 | 1234567890123345\n||||12345  | None\nAlpha Numerals|*^[a-zA-Z0-9\\]+$|Accepts both alpha characters and numbers from 0-9|johnjacob123 | johnjacob123\n||||johnjacob*&1  | None\nAccept Alpha Numerals with Special Characters|^[a-zA-Z0-9_-*/%&\\]+$|Accepts both alpha characters and numbers from 0-9 including special characters|johnwick@123 | johnwick@123\n Scrub first 4 characters in a string|^[\\s\\S\\]{0,4}|Selects only  first 4 characters of any string| DUNE_world |DUNE\n||||123456 | 1234\nScrub Last 3 characters in a string|.{3}$|The dot operator represents characters from the end, so number 3 denotes to scrub last 3 characters| DUNE_Rocks | cks\n||||123456 | 456\nScrub only first name from Full Name|^[^,-. \\]*|This Regex returns the first name that is separated by hyphen(-) or comma(,) or space| Alex, Feliciano |Alex\nScrub only last name from Full Name|(?<=[,-. ]).*|This Regex will returns the last name that is separated by hyphen(-) or comma(,) or space|Alex- Feliciano| Feliciano\nZIP code Validator|^\\d{5}[-\\s]?(?:\\d{4})?$|Accepts 9 digit zip code and can be separated by a hyphen (-)|12345-6789 | 12345-6789\n||||1234| None\nSSN Number Validator|^\\d{3}-\\d{2}-\\d{4}$| Accepts 9 digits SSN code that is divided into first 3 digits next 2 and last 4 digits separated by hyphen.|12345-6789 | 12345-6789\n||||1234| None\nAccept Valid Date|MM/DD/YYYY format - ^(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])\\/(19\\|20)\\\\d{2}$| The pattern  (0[1-9]\\|1[0,2]) represents 1 to 12 digits which is applicable for month validation. '|22/03/2003| 22/03/2003\n||DD/MM/YYYY format - ^(0?[1-9]\\|[12][0-9]\\|3[01])\\/(0?[1-9]\\|1[0-2])\\/(19\\|20)\\\\d{2}$|( 0[1-9]\\|[12][0-9]\\|3[01]) - This Regex represents numbers from 0 to 31 for date validation.|32/07/2005 | None\n||YYYY/MM/DD format - ^(19\\|20)\\\\d{2}\\/(0?[1-9]\\|1[0-2])\\/(0?[1-9]\\|[12][0-9]\\|3[01])$|(19\\|20)\\d{2} - This Regex accepts dates from 1900's and 2000's, with bar separates '/|2022/12/22|2022/12/22\n\n---\n**CHEAT - SHEET**\n|REGEX|DESCRIPTION|\n|---|---|\n|  .| Matches Any Character\n|\\d|  Digit (0–9)\n|\\D| Not a digit (0–9)\n| \\w | Word Character (a-z, A-Z, 0–9, _)\n| \\W| Not a word character\n| \\s| White space (space, tab, newline)\n| \\S| Not white space (space, tab, newline)\n| \\b| Word Boundary\n| \\B| Not a word boundary\n| ^| Beginning of a string\n $| End of a String\n [  ]| matches characters or brackets\n [^ ]| matches characters Not in brackets 14. | = Either Or\n ( )|  Group\n *|  0 or more\n +| 1 or more\n ?|  Yes or No\n {x}|  Exact Number\n{x, y}| Range of Numbers (Maximum, Minimum)|false|true|true|4|3.3 Commonly used Regular Expressions|82
761|TresataSupport||****\n\nLet's have a quick recap of the journey we had in Connect step. We started by understanding the significance of Connect, moved on to learn the screen controls, and finally went ahead to add our resolution logic to link data together.\n\nIn this post, we shall look into the criteria on which the selected fields are coming along together.\n\n**Configure Connector Type**\n\n![Connect_Configure_Connector_Type|690x359](upload://zQ0b057YFZOiOvP3Gs6ifZtgMXh.png)\n*Connect: 4.0*\n\nNow that canonical fields are added, and even created internal linkages by adding parentheses in required places, but on what condition are these fields getting linked together? In addition to connect when the field values are same, there are a few other ways in which values in two fields match for two records, some specific to certain types of fields.\nYes, here is the answer to it. Tresata offers different type of Connectors that decides how records will be linked. Here is the brief insight on all connector types.\n\n1. Same: This connector type converts strings into lowercase and creates a match when there is exact comparison. This matcher type doesn't consider *null* values.\n\n2. Name: The name matcher can be applied to only Name field. The main functionality of this is that it parses raw name string into firstName, lastName, middleName, middleInitial, nameTitle, suffix and performs matching on the parsed values.\n\n3. Address: This Address matcher works similar to Name Matcher, and can be applied only on address fields. This address matcher will accept the raw address string and parse that into house number, road, level, unit, city, postcode, state and country. Then continues to match values based on the parsed fields.\n\n4. CompanyName: Company Name Matcher can be applied to only Company Name. As the above matchers, this will parse raw company name string into Company name, activity, region, structure and legal. After parsing, it performs matching operation on the basis of these parsed field values.\n\nUsers can choose one of the Matcher type from the above mentioned options to match their records.\n\n**Initiate Connect**\n\n![Initiate_Connect|690x359](upload://cva8UWrwOUFHy66jZnJGq4v3ZhB.png)\n*Connect: 4.1*\n\nWe have successfully reached the final part of CONNECT. After choosing the right canonical fields and its corresponding  connector types we are all good to execute the logic. As shown in screen 4.2 click on Initiate Connect button to start the execution. Users can go back to make any changes to their logic anytime before clicking on this button.\n\nThis concludes the Connect Step. Execution could take place anywhere between 30 to 1 hour for a small dataset, sit back and relax for a bit until Tresata completes doing this magic resolution. Feel free to post any queries you may have about this step on Community.\n\nCheers..!!!|false|true|true|4|4.4 Executing Connect Step|85
760|TresataSupport||Now that all the elements of the Connect step have been explained, it's time to have a walk through configuration in connect step and dive deep into creating connection logic to link records together.\n\n**CREATE CONNECT CONFIGURATION**\n\nThe first step to configuring connect is identifying what type of step or combination of steps best suits the user's case. Details about the available types of steps can be found in this post, but to summarize:\n* *Resolve*: Each record within the selected sources can connect with all the other records included in the sources according to the logic specified in the resolve step. Each cluster of records that connect together here get a unique id that differentiates one cluster from another which is known as a **Tresata Id**.\n* *Against*: Directional linkage, it connects one or more records from the selected sources on the "From" directory to at most one from the "To" directory according to the logic specified in the against step. It is mostly used to link records from transactional sources to those in reference sources. These transactional records are also given the same Tresata Ids as the record from the reference source to which they are connecting.\n\nThe choice of the step type, is heavily dependent on the sources, the user plans to connect with that logic. If the user wants to connect on only reference sources, they will use the *resolve* step for that but if the user then additionally want to connect the transactional sources on the resolved reference sources, they can go with the *against* step and specify *"from"* as the transactional sources and *"to"* as the reference sources.  The end result the connect step will be generation of Tresata Ids that will uniquely identify an entity and consists of multiple records from different sources (reference and transactional), everything about that entity under a single Id.\n\n**Source Selection Process**\n\n In *screen 3.0* the source selection process is shown for a *resolve* step. \n\n***PRO TIP***: *Remember, the **against** step allows connecting many records from transactional sources (transactions, purchases, bookings) to at most one record from reference data sources (clients, customers, members) since each transaction is unique to a specific type of entity.*\n\n![Connect_Add_Data|690x359](upload://hhpIAkbt9c8W74XXMlPxHAP5Vvp.png)\n*Connect: 3.0*\n\nAs shown in *screen 3.0*, the user can select the required dataset by clicking on the **(+)** in the *"Add Data Sources"* section. Once clicked, it will present the list of available sources and allow for real-time filtering while typing the name of the one to be added. Without choosing at least one source for each category (one category for *resolve*, two for *against* - *from* and *to*) the rest of the configuration panel is in a disabled state.\n\n-------------------------------\n**Creating Connect Logic**\n\nUpon selecting data sources, the canonicals included to **at least one** of the selected sources gets enabled on the *Canonicals* right panel. The panel includes:\n\n* ***Selected Sources (#)***: The canonicals included in **at least one** of the selected sources for this step.\n* ***Others (#)***: The canonicals not included in any of the selected sources for this step.\n* ***Color Coded Indication***: Based on the population of the canonicals. If the canonical is included in multiple sources, it is color coded based on the average across all of them. It allows user to plan whether to include a canonical in the logic. In *screen 3.0* the source selection process is shown for a *resolve* step.\n\nHovering over the canonicals, the user is able to see the exact percentage populated for each source, which enables more efficient connection logic.\n\n***PRO TIP***: *Choosing highly populated fields for Connect logic, ensures that most of the records will have values for those fields and thus, will be eligible to be checked for connections. If the least populated fields are present in the connection logic, least connections will be created, as empty values result in records being excluded from the linking process.*\n\n\n![Connect_Analyse_Canonicals|690x359](upload://83cgTO7lGRsgNRvpyzw9pqgGFlf.png)\n*Connect: 3.1*\n\n--------------------------------------------------------------------\n\nNow, After the user has decided the step type and has seen what canonicals are available in the selected sources to configure connection logic for that step, what is left is actually identifying what combination(s) of fields, if matching, define two records as describing the same entity and thus, form a connection. \n\nThe CONNECT strategy is heavily related to each use case. For example, different fields are used define a unique person than those used for a unique company. On a high level:\n\n* ***Connecting people***: name, phone, email, ssn (or id, passport etc), address, state, city, country, brithdate, gender and more.\n* ***Companies***: name, address, state, city, country, classification, date_of_incorporation, tax_code and more. \n\nSo for the first case, *name+phone* can identify a unique individual and so does *name+email* or just *passport id*. In the second case, *name+address* can identify an individual company and so does *name+date_of_incorporation* or just *tax_code*. So there can be multiple such combinations which identify a unique entity. This is where the *Add Logic* option is used to add as any such combinations as possible to identify more and more connections. \n\nOf course this is not an exhaustive list but rather, an indication of some of the fields could be interesting for each use case. Permutations of those plus other fields not included in the list above might be enough to define that two records describe the same entity. But how does a user actually configures that logic? \n\nAs shown in *screen 3.2*, the user can drag and drop fields from the Canonicals to the specified area in the Add Resolution Logic panel. Each white box represents a combination that, if fully satisfied, will create a link between records. \n\n\n* **Add Fields to Resolve:**\n\n![Connect_Add_Fields_for_Resolution|690x359](upload://reqUw36JRiyaS9E5WLePMJ8Rn9t.png)\n*Connect: 3.2*\n\nAs we have left with only required fields for resolution, let's start to drag and drop the fields from Canonical List to Resolution Tab.\n\n* **Parentheses Action:**\n\n![Connect_Parentheses_Action:|690x359](upload://9LUfxDTDjqQp7y44x431m6a7l16.png)\n*Connect: 3.3.1*\n\n![Connect_Parentheses_Action:|690x359](upload://tmGGIC2k3aKmjYht55y1v33FI5m.png)\n*Connect: 3.3.2*\n\nAdding a Parentheses to a canonical field, creates an internal resolution. Screen 3.3.2, denotes that, a record link is created  only when of both address and city meet the threshold value that is set. This helps users to create multiple complex resolutions in just one step. There could be individual fields can also be used with fields within parentheses that leads to both internal and external resolution.\n\nThe above described steps shows an example of using Resolve method of resolution. Let's look into adding another step in the resolution process with Against method.\n\n* **Adding another Step of Resolution:**\n\n![Connect_Add_Step_2|690x359](upload://n1NsMePoy6de9X7GugpzVCsvpsC.jpeg)\n*Connect: 3.4*\n\nClick on the *Plus button* to add a new step as shown in the screen 3.4\n\n![Connect_Against_Method|690x359](upload://5SFlKf6MEyTIyFhMIkWk30RRhG6.jpeg)\n*Connect: 3.5*\n\nLet's choose Against Method of Resolution this time as an example. The steps to add fields shall remain same as we performed for Step-1. Drag and drop the required fields and their Target fields.\n\n\n---------------------------------------------------------------------\n* **Using Shields**\nAs explained in [4.2 Getting Started With Connect](https://community.tresata.com/t/4-2-getting-started-with-connect/544), *Shields* are essential to maintain integrity of connections and avoid forming incorrect links. They ensure that, regardless of whether connection logic is satisfied, if specific integrity safeguards are broken then links are removed between records. More specifically:\n\nShields operate across all steps, regardless of sources picked or logic defined. They include canonicals, that if inconsistent across records, connection **should not** be formed (birthdate: one person can't have two different birthdates, ssn: one person can't have two Social Security Numbers and more). While Connection Logic emphasizes on what **should** match, Shields define what **should not** match.\n\nA user should include in Shields fields that should be consistent and always the same for connected records (birthdates, ssn and more). If **any** of those fields is inconsistent, then the connection will not be formed. \n\n***PRO TIP***: *Remember, Shields operate on a higher level, across sources and steps. Thus, when defining them the user might be looking for a canonical that is not included in the sources picked for the current step. By clicking on *Others(#)* the user can find the rest of the canonicals and still use them as Shields in their configuration.*\n\n![Connect_Add_Shield_Fields|690x359](upload://1gPGxx3163fhX63ax3U1hiyKSKS.png)\n*Connect: 3.6*\n\nIf the user attempts to proceed to *Build Pipeline* without configuring any shields, a reminder is shown to highlight the importance of Shields to accurate connections as shown below.\n\n![Connect_Shield_Pop_Up|690x359](upload://vR64su0Nh4peUBSSkMnGlursxWS.jpeg)\n*Connect: 3.7*|false|true|true|4|4.3 Configure Connect Logic|85
759|TresataSupport||****\n\nIn the previous post, the importance of CONNECT for the process of gaining meaningful insights from user data is highlighted. But what are the main CONNECT configurations and how do they differ from each other? Answering the above is the main purpose of this post!\n\n**CONNECT**\n\nStarting from the top, first one notices the HeatMap, that can give meaningful insights as to what fields are populated & unique enough to contribute to accurate linkage.\n![Connect_HeatMap_Button|690x359](upload://dSmwoNDxURJhXdf4VB5tZtfDZCe.png)\n*Connect: 2.0*\n\n![Connect_HeatMap_View|690x359](upload://uVVBRPbd4aZQY37MX1eKxRFxt7d.png)\n*Connect: 2.1*\n\nAs shown in screen 2.0, click on the "View HeatMap" button to reach screen 2.1, including the HeatMap as generated in PROFILE. This way, the user can make informed decisions as to what fields will contribute the most to effective record connections.\n\n![Connect_Screen_Highlights|690x359](upload://raQZrBeLj5eh0FXUfpQ829kVIzd.jpeg)\n*Connect: 2.2*\n\nAs seen in screen 2.2, there are two standard methods in which users can create their logic to link the records together. They are:\n\n1.  **Resolve:**  This resolution type allows for any records within the selected sources to connect against any other records from the same and the rest of the selected sources according to the logic specified on the resolve step.\n\n* *For example, as seen in a previous post on [significance of connect](https://community.tresata.com/t/4-1-connect-its-significance/542), if user wants to know if Helen is the returning customer, they need to connect records' PII (name, address, birthdate and more) with past ticketing and booking purchases to identify whether she has purchased tickets in the past. Using  "**Resolve**" logic, they can match any record from the Ticketing source, to any other record from either Ticketing or Booking. If this matching process brings many records together, they can identify Helen as a returning customer.*\n\n2. **Against:** This resolution type, is a directional matching process. In detail, it attempts to connect records from a pool of source(s) (mentioned as "***from***") to at most on record of another pool of source(s) (mentioned as "***against***"). This step is particularly useful when connecting transactional data sources to reference ones (purchases to customers, transactions to clients and more). This is a many to one step, which means that since there can be multiple transactions corresponding to an entity, all these transactions can be attached to that same entity.\n\n* *After resolving all the booking and ticketing information together, there exists a common identifier for all the purchases Helen (or any customer for that matter) has with FunAirways. However, how to know whether those purchases are done by a member of their loyalty clients? They can attempt to connect all those records with one record on our Loyalty source (each record on the Loyalty source is unique, since each customer has a unique Customer_Loyalty_Number). Matching multiple transactions (bookings and ticketings) against client records is a classic example of an ***against*** resolution step.*\n\n3. **Steps:** CONNECT comprises of many steps, each one defining different ways to connect records for the selected sources within that step. Not all sources should connect with each other based on the same logic, look at the example above: Ticketing and Booking connected with each other with a resolve on PII information (canonicals like name, email, address and more). However, for Ticketing and Booking to connect to Loyalty (FunAirways loyal customers data source) the unique Customer_Loyalty_Number canonical is enough to bring them together with an against step. That flexibility is introduced to the user via steps.\n\n4. **Add Data Sources:** Prompts the user to add data sources to the selected step. Only the records from the selected data sources will be the only ones considered for matching with the configured logic within the step. \n\n5. **Canonicals:** Canonicals Tab is automatically populated immediately after the Data Source(s) is added. Those are the fields that can be used to build the logic for the step and define how should records for the selected sources connect. To further assist the process, upon hovering over the canonicals, the user can see how populated they are, which is an important indicator to how much each field can contribute to the connection process. \n\n6. **Add Resolution Logic:** That is the place where the connect logic is specified. As should in *screen 2.2*, there is a specified gray box where the user can drag and drop fields accordingly. Each box defines a combination of canonicals that, if matching, create a connection between two or more records. \n\n7. **Add Link SHIELDS:** In order to avoid incorrect connections, Tresata allows the user to define "shields", i.e. fields that if they have different values, the connection is incorrect and should be broken. \n\n* *Imagine a scenario where FunAirways reolves the list of passengers for one of their international flights with a list of people forbidden from entering that country. Now assume that for that logic, they use **name, email, phone, and citizenship**. According to that logic, one passenger, John Doe, seems to have connected with the list of **flagged** people and thus, should be denied during the boarding process. However, the manager of FunAirways, notices that the two records, while having similar PII (name, email, phone and citizenship) actually have different birthdate, idnicating that they are different people. Adding birthdate as a **SHIELD** would prevent that connection and improve the accuracy of the CONNECT step.*\n\n8. **Build Pipeline:** To proceed in CONNECT, the user has to first click on the "**Build Pipeline**"  button to enable Tresata's engine to calculate the pipeline for connections as defined by the user provided logic.\n\n\nWith this we have made ourselves comfortable with all the features Tresata provides for CONNECT phase. In our next post, lets see how to create our first resolution logic efficiently. Stay Tuned...!!!|false|true|true|4|4.2 Getting Started with Connect|85
757|TresataSupport||**SUMMARY**\n\nAfter the data has been cleaned and prepared, the next step is to identify and connect records across various data sources and soiled systems, so that the user has a more holistic view of a unique entity. \n\n*Seems simple, right? Not quite...*\n\nWhen dealing with multiple, diverse datasets, records may contain different attributes or have variations in how they represent the same entity. CONNECT allows the user to integrate these disparate pieces of information for each record into a more complete and accurate representation of the entire entity. \n\nBut why is this important and how does this help businesses grow? This post will aim to answer those two questions!\n\n**WHAT IS CONNECT**\n\nTo better understand the power of CONNECT, it may be easier to describe the problem using a real world example:\n\nHelen is a travel enthusiast always flying with the same airline company, FunAirways. Now, let's imagine each interaction Helen has with FunAirways as she books her upcoming flight to Greece. First, she books her round-trip ticket via the FunAirways website. Then, on the day of her flight, she checks in to her flight at the airport and purchases two checked bags at the counter. Next, she settles in to her flight and orders a smoothie from the flight attendant. Lastly, she arrives in Greece and heads to the rent-a-car counter, where she plans to pick up the car she reserved through FunAirways' website (using their trusted partner, FunCars, of course!). \n\nThat amounts to four separate interactions with FunAirways during her travel journey! What makes things difficult is that the records for each of those interactions are located in separate systems (i.e. the booking system is completely different than the in-flight services system). Thus, if FunAirways wanted to gain a comprehensive understanding of Helen, or any of its other customers, they would have a difficult time doing so. \n\nNow, let's make this problem even *more* difficult. Let's imagine that Helen used her home phone number and home address to book her ticket. However, the \n\nHow can FunAirways:\n\n* Identify that Helen is a returning customer, even though not a loyalty member, that constantly chooses them to fly with?\n* Identify patterns in Helen's behaviour to personalise their services (perhaps offering her a free smoothie during her next flight or even points for her next car rental)?\n\nCONNECT is Tresata's step for solving this problem. All different source come together, utilising a powerful entity resolution engine to identify unique entities within all the records, based on ML algorithms and user-defined logic.\n\n**WHY IS CONNECT IMPORTANT**\n\nBy creating a comprehensive, 360-degree view of each unique entity, CONNECT enables enterprises to understand an entity's characteristics, behaviors, and interactions across various contexts. This understanding allows businesses to enhance customer loyalty, operational efficiency, and make smarter decisions, achieving these goals faster than their competitors. This business model is employed by companies like Amazon, Google, and other FAANG members. These companies optimize every process and interaction by gaining deep, dynamic insights into individual customer behaviors and preferences. This approach facilitates the hyper-personalization of each customer relationship, which we, as consumers, have come to expect, thereby fostering unparalleled loyalty. By demonstrating to customers that they know, understand, and appreciate their unique preferences and behaviors, these companies ensure customers keep coming back.|false|true|true|4|4.1 Connect & its Significance|85
754|TresataSupport||**SUMMARY**\n\nAs we have established a functional workflow, the crucial next step is to monitor its progress and address any errors that may arise. This post outlines various methods to effectively check on the workflow.\n\n**USER ACTIONS**\n\n![Orchestrate_Progress Bar|690x359](upload://2Psgivq7Mtm4UANOvRZENnds1EB.png)\n*Orchestrate: 2.0*\n\n* *Progress Bar:*\n Users can choose just one stage of the workflow to all stages of the workflow. Based on the selected stages, user can view the progress of their running workflow as shown in the screen 2.0\n\n![Orchestrate_Restart_Workflow|690x359](upload://xyPwqtZ3wLI8gJexxTcdNI5FTy6.png)\n*Orchestrate: 2.1*\n\n![Orchestrate_Restart_Workflow_Approve|690x359](upload://decmLbKTaqzCNLdiDKUCSnxQJYw.png)\n*Orchestrate: 2.2*\n\n* *Restart Workflow:*\nWhen there is a change in workflow or rerun the workflow, users can easily do so by using the restart option as shown in the screen 2.1. After which there is a pop up on screen to confirm the restart option as seen in screen 2.2\n \n\n![Orchestrate_Cancel_Workflow|690x359](upload://rvaZ7ggh1kvt4F1Zh8mbUDYMp9r.png)\n*Orchestrate: 2.3*\n\n* *Cancel Workflow:*\n Users can just cancel the running workflow, if there is a situation that demands a change in the scheduled run.\n\n* *Start, Edit and Delete Methods*\n\n![Orchestrate_Start_Workflow690x359](upload://sdqEgZqYqGPutVqS3HyjtpO5XMb.png)\n*Orchestrate: 2.4*\n\n1. Start: Users can start the run whenever they prefer to irrespective of the scheduled time as shown in screen 2.4\n\n![Orchestrate_Edit_Workflow|690x359](upload://2g4cs8EM7ymGAqINH209cAyMJSX.png)\n*Orchestrate: 2.5*\n\n2. Edit: Users can edit the timelines by clicking on the “pencil button” to change duration, time etc to anything that is according to user requirements as seen in screen 2.5\n\n![Orchestrate_Delete_Workflow|690x359](upload://zpmENySIOJvrNrhvQ5xOwYKCOfQ.png)\n*Orchestrate: 2.6*\n\n3. Delete: Looks like user made a mistake while scheduling or chose a wrong workflow? Or user no longer want the schedule to happen ? Never mind, user can choose the workflow they just scheduled and click on delete option to remove them as shown in screen 2.6.\n\n**THINGS TO REMEMBER IN ORCHESTRATION**\n\nThere are few important points to remember while setting up the workflow to orchestrate\n\n* The name of the workflow can not be changed. Once chosen in the beginning shall be the same name to all of the scheduled runs too.\n*  The name of the workflow can not have any special characters or can not have duplicated names.\n* Scheduled workflow can be changed and deleted at any point of time.\n\nFinally this completes all stages in the workflow. We hope this journey was comfortable and smooth. Please feel free to post any queries that you could have in community and we will help you sort the issue..|false|true|true|4|7.2 Monitoring Orchestrated Workflow|83
753|TresataSupport||Managing time efficiently is the key for the fast paced world. If we could automate the workflow created once, that shall run automatically at selected time. Yes. Tresata offers users to run their workflow from profiling their data to having an enriched data in just one click. The steps to be followed to orchestrate workflow is  discussed in this post\n\n**ORCHESTRATE THE WORKFLOW**\n\nAfter creating a complete workflow end to end, users can now automate them to run by itself in the internal that is set.  First click on *Automate Workflow* button to get started with Orchestration\n\n![Orchestrate_Automate_Workflow|690x359](upload://84NhJJmQXya7AI0AxIj25DvBicC.png)\n*Orchestrate: 1.0*\n\nThere are two types of Orchestration Techniques, that is provided in product. One being Manual and the other being Automatic Orchestration. Let's look into them individually to know how to use it.\n\n* MANUAL ORCHESTRATION\n\n![Orchestrate_Manual_Method|690x359](upload://mVRX3zZdNTvEUZtiyoxNIle3Vu7.png)\n*Orchestrate: 1.1*\n\nThe screen above shows how Manual orchestration method looks like. Whenever user has a workflow ready to be scheduled, they can select the workflow required to run in using the search bar. The workflow can just run one step like profiling or two steps like Profile and Prepare or user can even have an end to end workflow inclusive of all steps from from profile to enrich.\n\nNow select the schedule type to be *Manual* and then clicking on *Confirm & Orchestrate* button will trigger the workflow run. Since it is Manual method, workflow is set to run only when user desires.\n\n* AUTOMATIC ORCHESTRATION\n\nUnlike manual method, automatic method of orchestration as the name suggests, it runs automatically at the selected time interval.\n\n![Orchestrate_Automatic_Method|690x359](upload://c6tFl0nUgjiWj7I70PtIBi7jBhH.png)\n*Orchestrate:1.2*\n\nSelecting Automatic method, will open another window as seen in the screen 1.2, that allows the user to choose interval with the simple drop down button. \n\n1. Duration - Here users can select the duration, it could be day, month or even year. The workflow kicks off automatically when that time is met\n2. Time - Users can set hours and minutes at which they want to execute the workflow.\n3. If users select daily at 1 pm est, the workflow is run without any human intervention everyday automatically\n4. User has to be sure to know the steps that they want to run automatically.\n\nJust like we confirmed in Manual method, go ahead and click on  *Confirm & Orchestrate* to trigger the workflow run. From this point, the workflow gets kicked off automatically when the set time is achieved.\n\nThe more information about monitoring the scheduled runs will discussed in the next posts...!! \nStay Tuned..!!|false|true|true|4|7.1 Workflow Orchestration|83
744|TresataSupport||**SUMMARY**\n\nOnce all raw fields have been tagged and canonical fields have been created, the user must start to think about how each field should be standardized. Given that each data source is different, it is likely that you will have various different canonical fields. Thus, your cleaning methods of these fields will inevitably vary (you would not want to clean the alphanumeric field, email, in the same way as a numeric field like a phone number). \n\nNow, you might be wondering...how will I know what cleaning should be applied to each field? Tresata to the rescue! Tresata offers users a wide range of cleaners that can easily be applied to remove outliers and inconsistent values. See below for a step by step walk through.\n\n**TYPES OF CLEANERS**\n\nThere are two standard types of cleaner that TRESATA offers as listen below.\n\n* **GLOBAL CLEANER**:\n\n![Prepare_Global_Cleaner|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 2.0*\n\n As the name suggests Global Cleaners are those that are applied to all the canonicals of all the data sources automatically in one click. SAM chat-bot suggests the global cleaners like Null cleaner and Trim_Lower in order to standardise data across all canonical fields.\n\n* **FILED SPECIFIC CLEANER**\n\n![Prepare_Individual_Cleaners |690x359](upload://AeZofRunEkAlQ1gxMZA75UkPox1.png)\n *Prepare: 2.1*\n\nTRESATA offers a wide variety of pre-built cleaners that can be applied to your canonical fields. To make the process even easier, our SAM suggests a few standard cleaners based on the kind of data that you're working with. These cleaners help to clean the raw data making sure that data with correct format moves to the next stages of TRESATA. In order to use SAM suggestions you can simply hit the "APPLY" button so that the selected cleaners will be applied automatically for the chosen canonical fields. \n\n**CUSTOM CLEAN YOUR FIELDS**\n\nFirst, choose the field that should be cleaned from the list of canonical fields on the left. \n\n![Prepare_Select_Canonical_Field|690x359](upload://b5NaZM0LYdi5YsoQw7DJdep0UlN.png)\n*Prepare: 2.2*\n\nFrom the list of available cleaners, select the most appropriate based on the nature of your canonical. \n\n**TIP:** Click on each cleaner for a brief description and example so that you have a better idea of how your field will be cleaned. \n\nOnce you decide on a cleaner, just click on, "Add Cleaner To Field" to apply it to the canonical.\n\n![Prepare_Add_Cleaner|690x359](upload://8WdkGOYhaD50zTb0pV35RQ0xMRu.jpeg)\n*Prepare: 2.3*\n\nIf you wish to edit the cleaner or add additional cleaners to the same field, simply use the "Edit" option as shown below. You can also view all the cleaners that were applied by clicking on the radio button "View Applied Cleaners" and check how the cleaners work together by providing a sample test string. Additionally, if a cleaner is no longer required, you are able to use this same option to delete the unwanted cleaner.\n\nEach time a cleaner is applied successfully, a notification will appear on the top of the screen. Once you feel happy about all the cleaned fields, you can click on "*Mark Complete*" so that you can move to the next data source for cleaning messy data.\n\n![Prepare_Edit_Cleaner|690x359](upload://6gN7qiS7DWDhZRe0LkamaaYelMD.jpeg)\n*Prepare: 2.4*\n\nAs you are going through this process, it is easy to lose track of the cleaners that have already been applied. Use the "View Applied Cleaners" button option present at the bottom of the screen for a quick glance of all cleaners that have been applied to a field. Additionally, use the "View Heatmap" button on the top left to get a view of your tagged fields across sources. When you are happy about the cleaners used, remember to click *Mark Complete* to make sure the cleaning has been completed for the selected Data source. \n\n![Prepare_View_All_Cleaners|690x359](upload://ot6FwWr1KpFV29qOFShYJnbLF7a.png)\n*Prepare: 2.5*\n\nCheck out the next post for an in-depth look at some of the more advanced cleaners Tresata has to offer!\n\nThe final step of Prepare is to click on *Initiate Data Preparation* to apply all the cleaning that you just selected.|false|true|true|4|3.2 Cleaner Actions|82
743|TresataSupport||**SUMMARY**\n\nAfter using TRESATA's profile engine to gain valuable insights (# of records, % populated, top values, and more), the next step is to leverage this intelligence to clean the data accordingly. Getting this step right is critical because uncleaned data can have serious repercussions on the accuracy and reliability of a data product - inaccurate values and inconsistencies can skew results, potentially leading to incorrect decisions. Additionally, valuable time and resources are spent manually correcting data quality issues and managing the data, rather than deriving valuable insights from it. \n\nBy cleaning and standardising the data, you enhance the accuracy of the record linkage process, promote data integrity, and create a solid foundation for future analyses and data products. This post is dedicated to learning more about the first step in cleaning up messy data: canonical fields.\n\n**CANONICAL FIELDS**\n\nCanonical fields refer to a set of standardised, commonly recognised fields used to represent specific attributes of the data. These canonical fields serve as fundamental elements to analyse data, create pipelines and derive valuable insights. They form a consistent and uniform representation of data across different sources, establishing a common language and structure for the profiled data (a common schema across all sources).\n\nFor example, let's say you have two sources (Table-1 and Table-2). \n\n* Table-1 contains the raw field name "*Full_Name*", representing customer names \n* Table-2 contains the raw field name "*Cust_Name*",  representing customer names\n\nSince both fields represent the same attribute, you would tag each field as ***name***, resulting in the creation of a single, universal canonical field called "name" (refer to the Profile step for further information on tagging). \n\n***Note:*** The tags you assigned in the Profile step are **automatically populated as canonical fields** during the Prepare step. \n\n---\n**GLOBAL CLEANERS**\n![Prepare_Global_Cleaner_By_SAM|690x359](upload://957p6RtKoFz3x9BeKlV6nnKhcyI.png)\n*Prepare: 1.0*\n\nIn Screen 1.0, you can see an example of the canonical list for the data source **boromir-gb-1**. The user has tagged over 10 fields that will be used in the following steps. Before cleaning the data, you can validate that these canonical fields are accurately tagged, and can add or delete new ones based on the specific use case. Once you have confirmed the canonical list is complete, they will dive deeper into field-level cleaning.\n\nThe next post is dedicated to explaining different data cleaning methods in TRESATA. Check it out for more detailed insights on how to standardise your data!|false|true|true|4|3.1 Prepare & its Significance|82
742|TresataSupport||Heatmap is the last part of Profiling stage. They are the visual representation of data patterns and relationship between different fields across multiple data sets that was profiled. HeatMap is created using different tags that were assigned by you, making it a one place destination to have complete view of your data.\n\n**REVIEW HEATMAP**\n\n![Profile_Review_Heatmap|690x359](upload://AgT9S5a7KMK3qkrLzpGv16DHxAg.png)\n*Profile: 5.0*\n\nWhen you have completed tagging their critical fields, you will get access to Heatmap.\nAs Heatmap is created based on the tags assigned, it is crucial to have at least one tagged filed before proceeding to Heatmap. \n\nAs shown in screen 5.0, clicking on Review Canonical Heatmap button will display the final heatmap.\n\n![Profile_Heatmap_view|690x359](upload://r7lBAyIsfGdyeONwK9bxI1lurmw.png)\n*Profile: 5.1*\n\nScreen 5.1 shows the resultant Heatmap that is created for the profiled data sets.\n* **List of Tags:** List of Tags tab shows all the tags that was assigned by you. The tags act as different categories and shows all the fields that was assigned the same tag. These tags are then considered as canonical filed names, which will be used for cleaning the field, creating pipelines etc. \n* **Sources:** In the screen 5.1 we see boromir-gb-1, ticket and sales being 3 different data sets. Each source is again broken down into 3 sub divisions like filed names, # of Uniques and % of populated.\n* **Field Names:** This is the raw names of the fields that was profiled.\n* **# of Uniques:** Shows the total count of unique values in the field. This details will help to identify the diversity of the data.\n* **% of Populated:** This column shows the cumulative percentage of the data that is populated in the column. The color gradients are used to encode values. \nMore populated values are represented in shades of green to show that these fields are fit to consider for next stages. Gradually it turns orange when we see 50% of population and color red denotes the values are critically low data population.\n\n**HEAT MAP ACTIONS**\n\n![Profile_Heatmap_Sort_Filter_action|690x359](upload://zNXq7Pi7LWZyUvEKD2tlgvN0n2K.png)\n*Profile: 5.2*\n\n* The Heatmap allows you to sort values according to the sources. As shown in screen 5.2, clicking on upward or downward arrows will sort the values in Heatmap according to the preference chosen.\n* Hide and un-hide sources by clicking on radio button that present next the source name. The heatmap updates itself with every new change made.\n* The lock button is used to make any data source to remain unchanged.  \n* Similar to the actions on source level, hide and un-hide options are available to field names, # of uniques and % of populated values. One click to change the heatmap according to requirement.\n* After making the changes, simply click on Apply button to update the heatmap.\n\n**HEATMAP HOVER ACTIONS**\n\n![Profile_Heatmap_Hover|690x359](upload://dl41Hz0rgOFDc8FHQq46CMHJMXJ.png)\n*Profile: 5.3*\n\nYou can hide any tags on the Heatmap by easily clicking on the eye button in front of every tag\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://4t4R6GtiaaZBsPwcCHVufkTTkiq.png)\n*Profile: 5.4*\n\nWhen hovered on the name of the field, you can view the Top values with the total percentage of that value present in the data.\n\n![Profile_Heatmap_Hover_FiledNames|690x359](upload://3TvfD7KnSbunMOVxKEErVLy1oWk.png)\n*Profile: 5.5*\n\nIn addition the details shown in screen 5.4, users can also view Top patterns of the field with the percentage of population for more understanding.\n\n![Profile_Heatmap_Hover_Population|690x359](upload://hiuETNWAQ1z0lvJrdxH63QU59eg.png)\n*Profile: 5.6*\n\nScreen 5.6 shows the action when hovered over the percentage of population column. This shows the details of the percentage used for color code\n\n**NEXT STEP**\nWhen you are happy about the over all heatmap, you will be able to export them to a csv in just one click for further reference of their holistic profiled data.\n\nThis brings us to the end of Profiling step. If you are experiencing any problems, reach out to our community team or post your quetsions here on [Tresata Support](https://community.tresata.com/c/tresata-product-support/94)|false|true|true|4|2.5 Profile Heatmap|80
736|TresataSupport||After a detailed investigation on different fields of the dataset, organising and categorising them is essential to start working on your data. In order to do that, TRESATA offers a special feature known as "Tags." These Tags are essentially keywords or labels that you can assign to critical fields, such as name, email, phone, ID, and more.\n\nWhen these Tags are assigned, they serve as canonical fields, enabling you to generate a comprehensive Heat-Map at the end of Profiling phase. Not only that, these tags become canonical fields, upon which the logic to connect datasets together created.\n\n**ADDING NEW TAG**\n\n![Profile_Add_New_Tag|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 4.0*\n\nAs shown on screen 4.0 above, to all the critical fields, you can easily add a new tag simply by clicking on the add button shown at the bottom of the screen\n\n![Profile_Save_Tag|690x359](upload://s0kYJ9fVB9oX8e84eEKnjFqky50.png)\n*Profile: 4.1*\n\nWhen you have finished adding a tag, clicking on save button will retain the tags that are assigned as shown in screen 4.1\n\n![Profile_Edit_Tag|690x359](upload://rPVijBKDbIAwdYMZDg8xnRUv22a.png)\n*Profile: 4.2*\n\n![Profile_Delete_Tag|690x359](upload://1Y9JH8QNhktHn57xbO6kclETseC.png)\n*Profile: 4.3*\n\nThe screen 1.1 shows that, the tags that are already assigned can be edited to a new tag at any point while doing the investigation of Fields. Similarly, as shown in screen 4.3, you can also remove the tags when found otherwise.\n\n**Best Practices To Add a Tag**\n\n![Profile_Tags_with_no_special_characters|690x359](upload://96JTaN0JPzU4YgjOhjklt6plRQK.png)\n*Profile 4.4*\n\n* **No Special Characters**: As shown in the screen 4.4, refrain using any symbols or special characters as tags, instead use more descriptive names \n\n* **Only One tag per Field**: Each field can have only one Tag assigned to it.|false|true|true|4|2.4 Add Tags to Fields|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78
717|TresataSupport||Looking at statistics on a source level is not granular enough to really understand what's in the data, identify data quality issues or even categorise fields to fit your need and requirements. To do all that, you will want to have the understanding of information on a field level, with overall statistics per field, visibility into actual values etc. All that an more, are available in TRESATA, enabling you to get a holistic understanding of the data.\n\n**LEFT SIDE PANEL**\n\n![Profile_field_landing_correct|690x359](upload://lmHNwJrR3e3fjwwEKULF45f4Uss.png)\n*Profile: 3.0*\n\nAs shown on screen 3.0 above, in order for you to investigate a source per field, you need to click on the expand button next to the source name on the left side navigation panel. Doing so, the source's view gets expanded, revealing all the fields included as well as a search bar to quickly search for a specific one. Notice that on the left side panel, around each field name there are some elements:\n\n* **Tags**: Under each name, there is a tag to categorise what this field is about. If there is no tag, that means the field hasn't been tagged yet (default state). You can learn more about this **crucial** tagging step ***here***. \n* **% Populated**: Represents the cumulative percentage of the data that is populated in the column. It gives an idea of the data's completeness. Notice that the values are color coded: the greener the color is, the more populated the field is. As the color is gradually approaching red, that mean there are more and more missing values.\n* **# of Uniques**: Shows the total count of unique fields present in the column. It helps identify the diversity or distinctiveness of the data.\n\nNOTE: You can use the sorting functionality next to the search bar to re-order the fields according to population and uniqueness, with flexibility on the order (ascending or descending).\n\nUsually, highly populated and unique fields are considered good to use later in the TRESATA processes. While that depends on the use case, it's always good to note down findings utilising the Notes functionality, as shown ***here***.\n\nWhile those metrics are good for high level field understanding, there still could be problems that you can't identify unless seeing the actual values within a field. Imagine a scenario where a phone company is testing their phone numbers and for that exercise, create ten thousand records with 0000-000-000.. the data would look complete but in reality, this is bad placeholder data. Or even a scenario where, user input on phone numbers doesn't specify format, and users end up putting their numbers like 1234-123-123 while other prefer 1234123123. To solve this problem, TRESATA allows you to go **even more granular** to the actual values within the fields. \n\n---\n**FIELD LEVEL INFORMATION**\n\nAs shown on screen 3.0, the middle panel reveals overview level statistics on the top bar and value based information on the rest of the middle panel. Often patterns or values can get very long which can cause truncation. Hovering over the truncated value will reveal the whole string, as in screen below:\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.1*\n\nLooking at the value based information, you can see:\n\n* **Top Values**: Provides the top values that are most frequently populated in the column. It helps identify common or frequently occurring data values. often, by looking at the top values, it is easy to identify placeholder or bad values (i.e. 1234567890 phone number).\n* **Top Patterns**: The top recurring patterns observed in the column's data. Investigating this gives visibility on whether data within a column has standardised format (23-02-1999 or 23/02/1999).\n* **Top Formats**: Displays the most commonly used data format in the column. It helps identify the dominant data format or structure present in the column. \n\nKnowing that there is a problem isn't that useful if you can't understand how big of a problem it really is. That's why next to each of those, you can see the actual percentage those values hold within the data. Additionally, you can in real-time filter those values out of your data to identify how that would affect the overall statistics of that field as shown below:\n\n![Profile_field_unselect|690x359](upload://7ogxSFdoZ4dXZiy2MFidb9BexkD.png)\n*Profile: 3.2*\n\n![Profile_Field_Level_Hover_Over|690x359](upload://ps8mVq8uxOL7ZHOEFMbedGv4eIF.png)\n*Profile: 3.3*\n\nInvestigating that middle panel is a **very important step for a successful TRESATA workflow**, especially when the field being investigated is a critical data element (name, email, phone, id and more). During this process you can identify Data Quality problems, trend and more.\n\n---\n\n**SAM : SIMPLE AUGMENTED MODE**\n\nTresata's very own chatbot SAM, suggests the you to take make effective choices with it's AI powered  suggestion. When you land on the profile page, SAM suggests the tags that are most important for your data source based on the resolution type on which the product was created.\n\n![Profile_SAM_Tag_Suggestion|690x359](upload://9xDFgMboaXm2ryPasCnxpRt7W8T.png)\n*Profile: 3.4*\n\nThe screen above is the representation on how SAM is suggesting most critical fields, where you can tag them from your raw data. Additionally, completely understanding the data is important for **tagging**, which is what powers the remaining TRESATA steps and will be explained ***[here](https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport)***.|false|true|true|4|2.3 Field Level Investigation|80
716|TresataSupport||The first step to understand your data.. is ensuring all of it is present to be investigated! TRESATA enables you to do that by showing Overview Statistics, as a whole or per source, as well as information to ensure that this is the latest and greatest of your data.\n\n**PROFILE LANDING STATISTICS**\n\n![Profile_Overview_Statistics|690x359, 100%](upload://m1TgdgmuOsMC0JByXs0Q1Bmsep0.png)\n*Profile: 2.0*\n\nAs you proceed from SOURCE to PROFILE, this is the landing screen showing the high level statistics of what has been processed so far by the PROFILE job. At this point, there are two possibilities:\n\n* All of your sources are successfully profiled and the left "Profiled Data Sources" reflects all of them.\n* Some of your data sources are profiled and for the rest, the job is still pending. The left side panel shows only the sources for which the job has been completed and the statistics reflect those sources accordingly.\n\nNotice that on the left side panel, nothing is selected. That way, Tresata's engine will sum up the available metrics to give you a high level idea of **everything** that has been processed so far, across all the completed sources. Available metrics:\n\n* Number of Sources (Tables)\n* Number of Records (Rounded Up)\n* Number of Fields (Columns) \n\nBy looking at those statistics, you can identify whether records have been dropped, tables have been skipped or even if there are fields that haven't been processed. However, those statistics become more interesting when looked on a source level.\n\n![Profile_Overview_Per_Source|690x359](upload://aPtmte89jjM7lFgPwg4vrrBHAdh.png)\n*Profile: 2.1*\n\nNotice that to get to that view, you have enabled the "Selected All" option on the left panel, meaning that the information on the right side will include all the completed sources statistics, per source. The elements included on the right tab now are:\n* **Number of Records**: Records (rows) for this source.\n* **Number of Columns**: Columns (fields) for this source.\n* **Path**: Location for this source on the cloud storage system (provides information about the directory or folder structure). For usability, the "Copy to Clipboard" functionality is present.\n* **Profiled On**: The last profile date for this source. For the early versions of TRESATA, this is to ensure that what you are looking at is the latest version of your data.\n\nTo enable you quickly navigate through the right side panel, an auto scroll option is available. By clicking on the top right drop-down, you can see a list of all your sources (the ones selected from the left panel) and decide which one they want to investigate.\n\nLooking at those statistics on a source level makes it easier to identify **if** anything is missing and **where** it is missing from. Once you identify that nothing is missing, you can proceed to have an even more granular investigation of the data, on a field level (checkout [this](https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport) post to learn more).|false|true|true|4|2.2 Profiled Overview Statistics|80
708|TresataSupport||PROFILE is a crucial step in the flow. In this post, we will identify:\n\n* **WHAT** is the PROFILE step\n* **WHY** is it important\n* **HOW** should it be interpreted\n\n**WHAT**\n\nProfiling refers to the process of analyzing and understanding data sources to extract valuable insights. It involves examining the structure and content of the data. More specifically:\n\n1. **Structure**: refers to high level information about your data (# of records & fields), as well as field names and types (numeric, string and more). \n2. **Content**: refers to the actual values included on those fields. PROFILE will provide information to the user in regards to the Top-Values, Patterns and Formats included, overall non-empty population, number of unique values and more, all on a field level. \n\n**WHY**\n\nEverything described above is key metrics, but why? Why is seeing and understanding those metrics crucial for downstream operations? \n\nGaining knowledge about values for fields with millions or billions of records is an extremely difficult task. Identifying problems in the data (test values, placeholder "bad" data, multiple formats), data completeness (non-null values for a field) as well as the unique values per field (is there duplication? how much?) are all findings that will drive decisions on PREPARE and CONNECT. Consider the following example:\n\n***SCENARIO**: An airline wants to test their new promotion system, where all loyal customers get an automated email with personalized template and offerings. In order to test that system, they create 10000 different records with the value "test" for customer_name field and "test@airline.com" for customer_email. Two months later, a Data Engineer is tasked to clean the sources for downstream usage, but how will he know about those test records among millions of data points?*\n\nFor the above scenario, running PROFILE workflow and looking at the Top Values & Top Patterns returned, you should identify that:\n\n* There is an unusual 4-letter pattern for full name\n* Among the top values for email, test@airline.com is there and needs to get cleaned\n\nWith that knowledge, they can now proceed to cleaning the data, enabling accuracy on later usage.\n\n**HOW**\n\nSo, WHAT is PROFILE and WHY is important has been established. But HOW to utilize PROFILE flow to maximize what you get from it?\n\nFor you, the most powerful way to use PROFILE output is:\n\n* Ensure all of your data is profiled using the overview numbers of # records and fields profiled across all sources.\n* Making sure you look through your fields for unusual patterns, placeholder values, irregularities on formats or low populated fields and not those down for each source on your notes (*"Notes" icon on top right of your screen*) in order to not lose those findings. \n* Making sure you check on the Tresata Suggested Tags for each field (when they are available) and either approve them, if they accurately reflect the field you are investigating, or create your own tag (*PRO TIP:* There are some pre-configured common tags at your disposal to use). tagging is **essential** for a successful workflow\n* Investigate and understand the PROFILE Heatmap view as it is critical for decision making on the rest of the steps.|false|true|true|4|2.1 Profile: What, Why & How|80
689|TresataSupport||**SUMMARY**\n\nAt this point, the user has validated their source is the one needed for this Data Product and no problems have been detected. Now, the only thing remaining is adding it and proceeding to PROFILE.\n\n**ADDING A SOURCE TO CART**\n\nTo add a source to the Cart, the user has to complete the whole journey of:\n\n* Choosing a format and checking the schema\n* Checking at least one field for the First 10 values\n\nOnce both those actions are done, the *"Add To Selected Data Sources"* button will be enabled for the user to use as shown below:\n\n![SOURCE-values-filled|690x359](upload://yVDGPF3Ijq4Se6rZSwTBAne5DUV.png)\n*Screen: 3.0*\n\nClicking on the *"Add To Selected Data Sources"* button, will reflect on the counter seen next to the "Continue to Profile", and the source boromir-gb-1 will be visible on that panel upon clocking on it as shown below:\n\n![SOURCE-CART-remove-one|690x359](upload://nqSAMWit9bHkEthtTlHqEp1aAC2.png)\n*Screen: 3.1*\n\nWhile in the cart, the user has the ability to perform specific actions:\n\n* **Individual removal**:\nIf the user click on the button as shown on screen 3.1, then they will see a pop up asking for confirmation for this action (screen 3.2). According to that action, the source will either be removed from the cart or will remain as initially selected.\n\n![SOURCE-remove-one-messages|690x359](upload://2KGxHAJZCIt0aQieVme7X5HDaa4.png)\n*Screen 3.2*\n\n* **Mass removal**:\nWhen the user click on the *Select All* check box besides *"Data Source(s)"*, a "*Remove Selected*" button appears, giving the option for the user to remove all the selected Data Sources. The user can adjust their selection by unselecting specific ones and then perform the action by clicking on that button. Screen 3.3 shows that view while screen 3.4 shows the confirmation pop up.\n\n![SOURCE-remove-all-button|690x359](upload://13djyuXo7jVqFW475ls6oEiNvPt.png)\n*Screen: 3.3*\n\n![SOURCE-remove-all-pop-up|690x359](upload://t72PAg0lgDNFcg0GLqYtDh1nQT.png)\n*Screen: 3.4*\n\n* **Continue to PROFILE**:\n\nWhen selecting this button, the user has finalized their selections and is ready to move to PROFILE. Once clicked, the user will get a confirmation pop up as shown in screen 3.5 and upon validating, they will be redirected to the Profile job monitoring panel where they can track the progress of the PROFILE job (screen 3.6).\n\n![SOURCE-proceed-profile|690x359](upload://q1brrm6kWlgdX8dfnMfrO4ylk0k.png)\n*Screen: 3.5* \n\n![PROFILE-job-status|690x359](upload://57wEWqhXD2JmsFd2KzcePHFPB2y.jpeg)\n*Screen: 3.6*\n\nThat concludes the SOURCE journey. If you are experiencing any problems sourcing problems, checkout the post dedicated to error on the SOURCE step in this category or reach out to the Community!|false|true|true|4|1.3 Add Source And Continue To Profile|79
688|TresataSupport||**SUMMARY**\n\nLooking at the file structure, it's easy to navigate and reach to a file, but how can the user ensure that they are using the correct file for their Data Product? Tresata enables that through:\n\n* Easy access to the source schema to verify the fields included\n* Easy access to the source first 10 records of user's file, to avoid corrupted files and give visibility on the actual values!\n\nBut how to do all that?\n\n**GET SOURCE SCHEMA**\n\nIn Tresata, the schema of a source will reveal the source's structure, i.e. the fields included in that source. Looking at the schema before In order to do that, the user has to navigate to the file they want to investigate by using the left side navigation panel or applying a direct search query using the whole path. Once the user has reached the desired, the screen should look like screen 2.0:\n\n![Sourcing-nested-expanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Screen: 2.0*\n\nNotice in the middle panel, the user is now prompted to choose the format their file has. A list of acceptable file formats will be available in the expand dropdown next to the *APPLY* button. The list of the available formats are:\n\n**Formats**: *parq*, *csv*, *csvu*, *bsv*, *bsvu*, *tldsv*, *tldsvu*, *casv*, *casvu*, *avro*, *json*, *orc*\n\nThe user can use the applicable to their source format as shown below:\n![SOURCE-schema-apply|690x359](upload://veh4chAvVcdqYPpcc37l8xOSdwS.png)\n*Screen: 2.1*\n\nOnce the format is applied, if correct (if not, checkout the dedicated post on errors in SOURCE), a list of the fields for that source will be available as shown on screen 2.2 below:\n\n![SOURCE-schema-fields|690x359](upload://9vSr2fssCAtpVWJGAaONfNutzCU.png)\n*Screen: 2.2*\n\n**NOTE**: If the source has multiple partitions, user can still run this on the parent folder and as long as all the partitions have the same format and schema, there should be no failures.\n\nThis is the first verification point, where the user can validate whether the source they are looking at actually has the fields needed for their Data Product. If yes, the next step is checking out the First 10 records for those fields...\n\n**GET FIRST TEN**\n\nNow the user knows the structure of the data, but what about the underlying values? What if the data is corrupted to if, for some reason, the whole file is empty? All those and more can be answered by simply looking at the first 10 record values for the selected fields.\n\nTo check out the data the user has to select the fields (up to 4 fields at one time) as shown in screen 2.3 below:\n\n![SOURCE-search-selection|690x359](upload://jjsu3MSNy7kQpIuyMa2PYWQTEFf.png)\n*Screen: 2.3*\n\nNotice that in the screen above, the user has utilised the available search box to quickly search and select the fields they are interested in exploring. Upon selecting the fields, the user can now *APPLY* the selection and the screen will look like this:\n\n![SOURCE-values-filled|690x359](upload://7zhEYcMbKpJT8iigkXCKTgX9Ysb.png)\n*Screen: 2.4*\n\nAt this point, the user can take multiple actions:\n\n* **Unselect a field**: will reorder the middle panel, putting the unselected field first after all the selected ones. The right side panel showcasing the values won't change until the *APPLY* button is clicked. The user can now pick another field(s).\n* **RESET**: will unselect all the selected fields, allowing the user to select new fields. The right side panel showcasing the values won't change until the *APPLY* button is clicked. \n* **Expand**: will expand the right side panel to provide more real estate for the values of the 4 fields selected. The screen of the view is shown below in screen 2.5.\n\n![SOURCE-values-expanded|690x359](upload://ddyPaynyQveShjQB9p4564tUW1D.png)\n*Screen: 2.5*\n\nAt this point, the user has all the necessary information to make a good choice whether this is one of the sources needed for this Data Product. In the next post, we will explore how to add a source to the Cart and the *Continue to Profile* flow.|false|true|true|4|1.2 Get Information About Your Source|79
687|TresataSupport||**SUMMARY**\n\nNavigating a directory structure is critical for anyone who interacts with files regularly. A directory structure, also known as a file system, is a hierarchical organization of folders and files that helps users manage and access data. Being able to effectively find and identify sources within a file system can lead to significant benefits in terms of efficiency and productivity. While the process might seem straightforward, it can become challenging as directory structures become more complex. \n\nTRESATA alleviates this complexity by providing an easy-to-use, flexible interface for users to quickly navigate through all levels of their file system.\n\nIn the following post we'll give a walk through of how TRESATA enables the user to:\n\n* View all objects (folders and files) existing on a user's back-end\n* Navigate quickly through a given file structure \n* Search a directory for a file path\n* Star important files and selectively access them\n\n\n**VIEW FILE SYSTEM**\n\n![Landing-Sourcing|690x360](upload://at20ZiFZOBnKMX7VuMuU4qynGr2.png)\n*Sourcing: 1.0*\n\nLooking at Screen 1.0, user will see an overview of the their files system. The left side panel mirrors the object structure existing on the back-end, giving visibility to the user on what folders and files exist on their system. In this example, the user has six directories: *"usecases"*, *"tresata-generated"*, *"user"*, *"ascii-directory"*, *"tmp"* and *"demos"*.  \n\nFurther breaking down the left side *"Objects"* panel:\n\n1. Each table is a file that can't include more files nested inside, while a directory is a folder including other directories or files within it.\n2. Each directory will have an *expand* indicator on the top right of it box, which when clicked will reveal the nested folder and tables (see example below in Screen 1.1)\n\n**NAVIGATE FILE SYSTEM**\n\nOnce the user is familiar with their file structure, the next step is to move in to a specific directory so that they can view its contents and easily find the file they are interested in. \n\n![SOURCE-no-sources-added|690x361](upload://k0dJvVr7T6nf7gJpkCYwOAlUQ9E.png)\n![SOURCE-no-sources-added|690x359](upload://pbtOycwsOtSGzHhua11JxVGUt65.png)\n*Sourcing: 1.1*\n\nIn Screen 1.1, we can see that *usecases* has been expanded to reveal the directories nested within. Notice that there is a search box where the user can search for a specific file or directory and see the results returned in real-time. However, if the user does not know the exact name of the file they are looking for, they can continue to navigate through the available objects until they reach the specified file. \n\n![Sourcing-nested-epanded-final|690x362](upload://fleCAkjW9HCGbUHJlrw8FFQZUro.png)\n![Sourcing-nested-epanded-final|690x359](upload://tl2d4euShoojjeRYhU7CVcHHGSr.png)\n*Sourcing: 1.2*\n\n*Tip:* To return to the structure where *usecases* is shown as the parent directory, the user has to click to "**Go to usecases**" and the subdirectories under *usecases* will be displayed.\n\nGiven the complexity of a file structure, it is critical for the user to know the exact location of file so that they can return to it with ease. TRESATA automatically displays the location of their file as the user navigates further down the nested structure. Screen 1.3 shows a clear example of this. Notice that the path is hyperlinked - clicking on any of the directories there will filter the left side panel and render the nested folders/files within that directory. \n\n![SOURCE-truncated|690x359](upload://mxzd5MtHwTDb87PFDa4oPMqFXQh.png)\n*Sourcing: 1.3*\n\nAside from redirecting to a specific directory through the path, the user can also copy to clipboard by clicking on the button next to it as shown on screen 1.4.\n\n![Source-clipboard|690x359](upload://g3p0j7NbWxIQkwvCavvSuDUGVw9.png)\n*Sourcing: 1.4*\n\n\n**ADVANCED SEARCH**\n\nTRESATA has a universal search box with a "Search using file path" message. The user can paste a file path which, enabling a direct search that will be reflected on the left side *Objects* panel.\n\n**NOTE**: This is just the beginning. TRESATA's advanced search capabilities for SOURCE will be enhanced on new releases, allowing for many more ways for the users to directly search for their sources.\n\n**STAR RELEVANT FILES / DIRECTORIES** \n\nUsers may often need to access the same set of files or directories repeatedly, making it cumbersome to navigate through a complex file system each time to locate and apply transformations to those files. To simplify this process, TRESATA offers a feature that allows users to star files. Once starred, these files can be viewed separately, saving time and effort.\n\nTo star a file or directory, locate the desired file or folder and click on the star symbol located just before its name. When clicked, the star will turn blue as shown in screen 1.5.\n\nNow for displaying only starred files, click on the toggle next to *"Objects"* that has "Show Starred only" written beside it as shown on screen 1.6.|false|true|true|4|1.1 Navigate & Select Your Source|79
683|TresataSupport||This section contains the documents on the Profile step of the TRESATA. \n\n* https://community.tresata.com/t/2-1-profile-what-why-how/498?u=tresatasupport\n* https://community.tresata.com/t/2-2-profiled-overview-statistics/503?u=tresatasupport\n* https://community.tresata.com/t/2-3-field-level-investigation/504?u=tresatasupport\n* https://community.tresata.com/t/2-4-add-tags-to-fields/521?u=tresatasupport\n* https://community.tresata.com/t/2-5-profile-heatmap/527?u=tresatasupport\n* https://community.tresata.com/t/profile-full-walkthrough/669?u=tresatasupport|false|true|true|4|About the Profile category|80
682|TresataSupport||This category consists of all the relevant documentation that is required to complete the *"Source"* step in the process of creating a data product. This includes:\n\n1.1 Navigate & Select Your Source\n&nbsp;&nbsp;1.1.1 View all objects (folders and files) existing on a user’s back-end\n&nbsp;&nbsp;1.1.2 Navigate quickly through a given file structure\n&nbsp;&nbsp;1.1.3 Search a directory for a file path\n&nbsp;&nbsp;1.1.4 Star important files and selectively access them\n\n1.2 Get Information About Your Source\n&nbsp;&nbsp;1.2.1 Get Source Schema\n&nbsp;&nbsp;1.2.2 Get First Ten Records\n\n1.3 Add Source And Continue To Profile|false|true|true|4|About the Source category|79
681|TresataSupport||(Replace this first paragraph with a brief description of your new category. This guidance will appear in the category selection area, so try to keep it below 200 characters.)\n\nUse the following paragraphs for a longer description, or to establish category guidelines or rules:\n\n- Why should people use this category? What is it for?\n\n- How exactly is this different than the other categories we already have?\n\n- What should topics in this category generally contain?\n\n- Do we need this category? Can we merge with another category, or subcategory?\n|false|true|true|4|About the Tresata category|78


298|TresataSupport||<a name="civilized"></a>\n\n## [This is a Civilized Place for Public Discussion](#civilized)\n\nPlease treat this discussion forum with the same respect you would a public park. We, too, are a shared community resource &mdash; a place to share skills, knowledge and interests through ongoing conversation.\n\nThese are not hard and fast rules. They are guidelines to aid the human judgment of our community and keep this a kind, friendly place for civilized public discourse.\n\n<a name="improve"></a>\n\n## [Improve the Discussion](#improve)\n\nHelp us make this a great place for discussion by always adding something positive to the discussion, however small. If you are not sure your post adds to the conversation, think over what you want to say and try again later.\n\nOne way to improve the discussion is by discovering ones that are already happening. Spend time browsing the topics here before replying or starting your own, and you’ll have a better chance of meeting others who share your interests.\n\nThe topics discussed here matter to us, and we want you to act as if they matter to you, too. Be respectful of the topics and the people discussing them, even if you disagree with some of what is being said.\n\n<a name="agreeable"></a>\n\n## [Be Agreeable, Even When You Disagree](#agreeable)\n\nYou may wish to respond by disagreeing. That’s fine. But remember to _criticize ideas, not people_. Please avoid:\n\n* Name-calling\n* Ad hominem attacks\n* Responding to a post’s tone instead of its actual content\n* Knee-jerk contradiction\n\nInstead, provide thoughtful insights that improve the conversation.\n\n<a name="participate"></a>\n\n## [Your Participation Counts](#participate)\n\nThe conversations we have here set the tone for every new arrival. Help us influence the future of this community by choosing to engage in discussions that make this forum an interesting place to be &mdash; and avoiding those that do not.\n\nDiscourse provides tools that enable the community to collectively identify the best (and worst) contributions: bookmarks, likes, flags, replies, edits, watching, muting and so forth. Use these tools to improve your own experience, and everyone else’s, too.\n\nLet’s leave our community better than we found it.\n\n<a name="flag-problems"></a>\n\n## [If You See a Problem, Flag It](#flag-problems)\n\nModerators have special authority; they are responsible for this forum. But so are you. With your help, moderators can be community facilitators, not just janitors or police.\n\nWhen you see bad behavior, don’t reply. Replying encourages bad behavior by acknowledging it, consumes your energy, and wastes everyone’s time. _Just flag it_. If enough flags accrue, action will be taken, either automatically or by moderator intervention.\n\nIn order to maintain our community, moderators reserve the right to remove any content and any user account for any reason at any time. Moderators do not preview new posts; the moderators and site operators take no responsibility for any content posted by the community.\n\n<a name="be-civil"></a>\n\n## [Always Be Civil](#be-civil)\n\nNothing sabotages a healthy conversation like rudeness:\n\n* Be civil. Don’t post anything that a reasonable person would consider offensive, abusive, or hate speech.\n* Keep it clean. Don’t post anything obscene or sexually explicit.\n* Respect each other. Don’t harass or grief anyone, impersonate people, or expose their private information.\n* Respect our forum. Don’t post spam or otherwise vandalize the forum.\n\nThese are not concrete terms with precise definitions &mdash; avoid even the _appearance_ of any of these things. If you’re unsure, ask yourself how you would feel if your post was featured on the front page of a major news site.\n\nThis is a public forum, and search engines index these discussions. Keep the language, links, and images safe for family and friends.\n\n<a name="keep-tidy"></a>\n\n## [Keep It Tidy](#keep-tidy)\n\nMake the effort to put things in the right place, so that we can spend more time discussing and less cleaning up. So:\n\n* Don’t start a topic in the wrong category; please read the category definitions.\n* Don’t cross-post the same thing in multiple topics.\n* Don’t post no-content replies.\n* Don’t divert a topic by changing it midstream.\n* Don’t sign your posts &mdash; every post has your profile information attached to it.\n\nRather than posting “+1” or “Agreed”, use the Like button. Rather than taking an existing topic in a radically different direction, use Reply as a Linked Topic.\n\n<a name="stealing"></a>\n\n## [Post Only Your Own Stuff](#stealing)\n\nYou may not post anything digital that belongs to someone else without permission. You may not post descriptions of, links to, or methods for stealing someone’s intellectual property (software, video, audio, images), or for breaking any other law.\n\n<a name="power"></a>\n\n## [Powered by You](#power)\n\nThis site is operated by your [friendly local staff](/about) and *you*, the community. If you have any further questions about how things should work here, open a new topic in the [site feedback category](/c/site-feedback) and let’s discuss! If there’s a critical or urgent issue that can’t be handled by a meta topic or flag, contact us via the [staff page](/about).\n\n<a name="tos"></a>\n\n## [Terms of Service](#tos)\n\nYes, legalese is boring, but we must protect ourselves &ndash; and by extension, you and your data &ndash; against unfriendly folks. We have a [Terms of Service](/tos) describing your (and our) behavior and rights related to content, privacy, and laws. To use this service, you must agree to abide by our [TOS](/tos).|false|true|true|4|GUIDELINES|33
278|TresataSupport||Community is the heart of Tresata. Community guidelines are a crucial aspect of any online platform or community.  To ensure a respectful and safe environment for all Tresata Community Members, we have set the following guidelines:\n\n* Engage respectfully, professionally, and with integrity at all times\n* Describe the situation & context, not specific details\n* Never share sensitive or revealing information (related to people, products, or clients)\n* Keep informal conversations outside of the community\n* Use Tresata Community for all technical topics/ threads\n* When responding to a post, attempt to solve or progress the conversation productively\n* Search for duplicates before posting\n* Use proper grammar and spelling\n* Facts > opinions, post thoughtfully\n* If you think something contributes to the conversation or is the right answer, upvote it and vice-versa\n* Zero-tolerance for inappropriate, hurtful, or negative content\n* [Reminder] - This is an open community so these guidelines apply to both internal & external user engagement, act accordingly|false|true|true|4|Community Standards and Guidelines|4
245|TresataSupport||Welcome and congratulations on becoming a member of the **Tresata community!** \n\nTresata Community aims to provide a robust platform, where you can find everything about Tresata products, Industry Best Practices and a common forum to Exchange Ideas and Information. This interactive platform provides a self-serve engagement forum where you can go through various informative topics, provide comments, communicate with Tresata experts using Personal Chat options or Emails, etc. \n\nYou will find like minded, Technology Enthusiasts, Data Champions, Tresata Product Experts, and Subject Matter Experts on this Tresata Community. \n\nKnow about using the portal here:\n![image|690x329](upload://n72U8QITc9VRqqzBs68ZRcAgwT5.png)\n\n\n\n\n\n\nYou will see personalised cards displayed on the [landing page](https://community.tresata.com/) covering multiple topic categories with relevant posts, specifically for you. The **GET STARTED** section will help you use the downloaded product easily.\n\nYou can leverage the robust **Search** functionality to find topic you are interested and leave comments, vote for the topic, or even create a new topic if needed.\n\nFor any support required, do reach out to support@tresata.com|false|true|true|4|Welcome to Tresata Community!|4
298|TresataSupport||<a name="civilized"></a>\n\n## [This is a Civilized Place for Public Discussion](#civilized)\n\nPlease treat this discussion forum with the same respect you would a public park. We, too, are a shared community resource &mdash; a place to share skills, knowledge and interests through ongoing conversation.\n\nThese are not hard and fast rules. They are guidelines to aid the human judgment of our community and keep this a kind, friendly place for civilized public discourse.\n\n<a name="improve"></a>\n\n## [Improve the Discussion](#improve)\n\nHelp us make this a great place for discussion by always adding something positive to the discussion, however small. If you are not sure your post adds to the conversation, think over what you want to say and try again later.\n\nOne way to improve the discussion is by discovering ones that are already happening. Spend time browsing the topics here before replying or starting your own, and you’ll have a better chance of meeting others who share your interests.\n\nThe topics discussed here matter to us, and we want you to act as if they matter to you, too. Be respectful of the topics and the people discussing them, even if you disagree with some of what is being said.\n\n<a name="agreeable"></a>\n\n## [Be Agreeable, Even When You Disagree](#agreeable)\n\nYou may wish to respond by disagreeing. That’s fine. But remember to _criticize ideas, not people_. Please avoid:\n\n* Name-calling\n* Ad hominem attacks\n* Responding to a post’s tone instead of its actual content\n* Knee-jerk contradiction\n\nInstead, provide thoughtful insights that improve the conversation.\n\n<a name="participate"></a>\n\n## [Your Participation Counts](#participate)\n\nThe conversations we have here set the tone for every new arrival. Help us influence the future of this community by choosing to engage in discussions that make this forum an interesting place to be &mdash; and avoiding those that do not.\n\nDiscourse provides tools that enable the community to collectively identify the best (and worst) contributions: bookmarks, likes, flags, replies, edits, watching, muting and so forth. Use these tools to improve your own experience, and everyone else’s, too.\n\nLet’s leave our community better than we found it.\n\n<a name="flag-problems"></a>\n\n## [If You See a Problem, Flag It](#flag-problems)\n\nModerators have special authority; they are responsible for this forum. But so are you. With your help, moderators can be community facilitators, not just janitors or police.\n\nWhen you see bad behavior, don’t reply. Replying encourages bad behavior by acknowledging it, consumes your energy, and wastes everyone’s time. _Just flag it_. If enough flags accrue, action will be taken, either automatically or by moderator intervention.\n\nIn order to maintain our community, moderators reserve the right to remove any content and any user account for any reason at any time. Moderators do not preview new posts; the moderators and site operators take no responsibility for any content posted by the community.\n\n<a name="be-civil"></a>\n\n## [Always Be Civil](#be-civil)\n\nNothing sabotages a healthy conversation like rudeness:\n\n* Be civil. Don’t post anything that a reasonable person would consider offensive, abusive, or hate speech.\n* Keep it clean. Don’t post anything obscene or sexually explicit.\n* Respect each other. Don’t harass or grief anyone, impersonate people, or expose their private information.\n* Respect our forum. Don’t post spam or otherwise vandalize the forum.\n\nThese are not concrete terms with precise definitions &mdash; avoid even the _appearance_ of any of these things. If you’re unsure, ask yourself how you would feel if your post was featured on the front page of a major news site.\n\nThis is a public forum, and search engines index these discussions. Keep the language, links, and images safe for family and friends.\n\n<a name="keep-tidy"></a>\n\n## [Keep It Tidy](#keep-tidy)\n\nMake the effort to put things in the right place, so that we can spend more time discussing and less cleaning up. So:\n\n* Don’t start a topic in the wrong category; please read the category definitions.\n* Don’t cross-post the same thing in multiple topics.\n* Don’t post no-content replies.\n* Don’t divert a topic by changing it midstream.\n* Don’t sign your posts &mdash; every post has your profile information attached to it.\n\nRather than posting “+1” or “Agreed”, use the Like button. Rather than taking an existing topic in a radically different direction, use Reply as a Linked Topic.\n\n<a name="stealing"></a>\n\n## [Post Only Your Own Stuff](#stealing)\n\nYou may not post anything digital that belongs to someone else without permission. You may not post descriptions of, links to, or methods for stealing someone’s intellectual property (software, video, audio, images), or for breaking any other law.\n\n<a name="power"></a>\n\n## [Powered by You](#power)\n\nThis site is operated by your [friendly local staff](/about) and *you*, the community. If you have any further questions about how things should work here, open a new topic in the [site feedback category](/c/site-feedback) and let’s discuss! If there’s a critical or urgent issue that can’t be handled by a meta topic or flag, contact us via the [staff page](/about).\n\n<a name="tos"></a>\n\n## [Terms of Service](#tos)\n\nYes, legalese is boring, but we must protect ourselves &ndash; and by extension, you and your data &ndash; against unfriendly folks. We have a [Terms of Service](/tos) describing your (and our) behavior and rights related to content, privacy, and laws. To use this service, you must agree to abide by our [TOS](/tos).|false|true|true|4|GUIDELINES|33
278|TresataSupport||Community is the heart of Tresata. Community guidelines are a crucial aspect of any online platform or community.  To ensure a respectful and safe environment for all Tresata Community Members, we have set the following guidelines:\n\n* Engage respectfully, professionally, and with integrity at all times\n* Describe the situation & context, not specific details\n* Never share sensitive or revealing information (related to people, products, or clients)\n* Keep informal conversations outside of the community\n* Use Tresata Community for all technical topics/ threads\n* When responding to a post, attempt to solve or progress the conversation productively\n* Search for duplicates before posting\n* Use proper grammar and spelling\n* Facts > opinions, post thoughtfully\n* If you think something contributes to the conversation or is the right answer, upvote it and vice-versa\n* Zero-tolerance for inappropriate, hurtful, or negative content\n* [Reminder] - This is an open community so these guidelines apply to both internal & external user engagement, act accordingly|false|true|true|4|Community Standards and Guidelines|4
245|TresataSupport||Welcome and congratulations on becoming a member of the **Tresata community!** \n\nTresata Community aims to provide a robust platform, where you can find everything about Tresata products, Industry Best Practices and a common forum to Exchange Ideas and Information. This interactive platform provides a self-serve engagement forum where you can go through various informative topics, provide comments, communicate with Tresata experts using Personal Chat options or Emails, etc. \n\nYou will find like minded, Technology Enthusiasts, Data Champions, Tresata Product Experts, and Subject Matter Experts on this Tresata Community. \n\nKnow about using the portal here:\n![image|690x329](upload://n72U8QITc9VRqqzBs68ZRcAgwT5.png)\n\n\n\n\n\n\nYou will see personalised cards displayed on the [landing page](https://community.tresata.com/) covering multiple topic categories with relevant posts, specifically for you. The **GET STARTED** section will help you use the downloaded product easily.\n\nYou can leverage the robust **Search** functionality to find topic you are interested and leave comments, vote for the topic, or even create a new topic if needed.\n\nFor any support required, do reach out to support@tresata.com|false|true|true|4|Welcome to Tresata Community!|4
298|TresataSupport||<a name="civilized"></a>\n\n## [This is a Civilized Place for Public Discussion](#civilized)\n\nPlease treat this discussion forum with the same respect you would a public park. We, too, are a shared community resource &mdash; a place to share skills, knowledge and interests through ongoing conversation.\n\nThese are not hard and fast rules. They are guidelines to aid the human judgment of our community and keep this a kind, friendly place for civilized public discourse.\n\n<a name="improve"></a>\n\n## [Improve the Discussion](#improve)\n\nHelp us make this a great place for discussion by always adding something positive to the discussion, however small. If you are not sure your post adds to the conversation, think over what you want to say and try again later.\n\nOne way to improve the discussion is by discovering ones that are already happening. Spend time browsing the topics here before replying or starting your own, and you’ll have a better chance of meeting others who share your interests.\n\nThe topics discussed here matter to us, and we want you to act as if they matter to you, too. Be respectful of the topics and the people discussing them, even if you disagree with some of what is being said.\n\n<a name="agreeable"></a>\n\n## [Be Agreeable, Even When You Disagree](#agreeable)\n\nYou may wish to respond by disagreeing. That’s fine. But remember to _criticize ideas, not people_. Please avoid:\n\n* Name-calling\n* Ad hominem attacks\n* Responding to a post’s tone instead of its actual content\n* Knee-jerk contradiction\n\nInstead, provide thoughtful insights that improve the conversation.\n\n<a name="participate"></a>\n\n## [Your Participation Counts](#participate)\n\nThe conversations we have here set the tone for every new arrival. Help us influence the future of this community by choosing to engage in discussions that make this forum an interesting place to be &mdash; and avoiding those that do not.\n\nDiscourse provides tools that enable the community to collectively identify the best (and worst) contributions: bookmarks, likes, flags, replies, edits, watching, muting and so forth. Use these tools to improve your own experience, and everyone else’s, too.\n\nLet’s leave our community better than we found it.\n\n<a name="flag-problems"></a>\n\n## [If You See a Problem, Flag It](#flag-problems)\n\nModerators have special authority; they are responsible for this forum. But so are you. With your help, moderators can be community facilitators, not just janitors or police.\n\nWhen you see bad behavior, don’t reply. Replying encourages bad behavior by acknowledging it, consumes your energy, and wastes everyone’s time. _Just flag it_. If enough flags accrue, action will be taken, either automatically or by moderator intervention.\n\nIn order to maintain our community, moderators reserve the right to remove any content and any user account for any reason at any time. Moderators do not preview new posts; the moderators and site operators take no responsibility for any content posted by the community.\n\n<a name="be-civil"></a>\n\n## [Always Be Civil](#be-civil)\n\nNothing sabotages a healthy conversation like rudeness:\n\n* Be civil. Don’t post anything that a reasonable person would consider offensive, abusive, or hate speech.\n* Keep it clean. Don’t post anything obscene or sexually explicit.\n* Respect each other. Don’t harass or grief anyone, impersonate people, or expose their private information.\n* Respect our forum. Don’t post spam or otherwise vandalize the forum.\n\nThese are not concrete terms with precise definitions &mdash; avoid even the _appearance_ of any of these things. If you’re unsure, ask yourself how you would feel if your post was featured on the front page of a major news site.\n\nThis is a public forum, and search engines index these discussions. Keep the language, links, and images safe for family and friends.\n\n<a name="keep-tidy"></a>\n\n## [Keep It Tidy](#keep-tidy)\n\nMake the effort to put things in the right place, so that we can spend more time discussing and less cleaning up. So:\n\n* Don’t start a topic in the wrong category; please read the category definitions.\n* Don’t cross-post the same thing in multiple topics.\n* Don’t post no-content replies.\n* Don’t divert a topic by changing it midstream.\n* Don’t sign your posts &mdash; every post has your profile information attached to it.\n\nRather than posting “+1” or “Agreed”, use the Like button. Rather than taking an existing topic in a radically different direction, use Reply as a Linked Topic.\n\n<a name="stealing"></a>\n\n## [Post Only Your Own Stuff](#stealing)\n\nYou may not post anything digital that belongs to someone else without permission. You may not post descriptions of, links to, or methods for stealing someone’s intellectual property (software, video, audio, images), or for breaking any other law.\n\n<a name="power"></a>\n\n## [Powered by You](#power)\n\nThis site is operated by your [friendly local staff](/about) and *you*, the community. If you have any further questions about how things should work here, open a new topic in the [site feedback category](/c/site-feedback) and let’s discuss! If there’s a critical or urgent issue that can’t be handled by a meta topic or flag, contact us via the [staff page](/about).\n\n<a name="tos"></a>\n\n## [Terms of Service](#tos)\n\nYes, legalese is boring, but we must protect ourselves &ndash; and by extension, you and your data &ndash; against unfriendly folks. We have a [Terms of Service](/tos) describing your (and our) behavior and rights related to content, privacy, and laws. To use this service, you must agree to abide by our [TOS](/tos).|false|true|true|4|GUIDELINES|33
278|TresataSupport||Community is the heart of Tresata. Community guidelines are a crucial aspect of any online platform or community.  To ensure a respectful and safe environment for all Tresata Community Members, we have set the following guidelines:\n\n* Engage respectfully, professionally, and with integrity at all times\n* Describe the situation & context, not specific details\n* Never share sensitive or revealing information (related to people, products, or clients)\n* Keep informal conversations outside of the community\n* Use Tresata Community for all technical topics/ threads\n* When responding to a post, attempt to solve or progress the conversation productively\n* Search for duplicates before posting\n* Use proper grammar and spelling\n* Facts > opinions, post thoughtfully\n* If you think something contributes to the conversation or is the right answer, upvote it and vice-versa\n* Zero-tolerance for inappropriate, hurtful, or negative content\n* [Reminder] - This is an open community so these guidelines apply to both internal & external user engagement, act accordingly|false|true|true|4|Community Standards and Guidelines|4
245|TresataSupport||Welcome and congratulations on becoming a member of the **Tresata community!** \n\nTresata Community aims to provide a robust platform, where you can find everything about Tresata products, Industry Best Practices and a common forum to Exchange Ideas and Information. This interactive platform provides a self-serve engagement forum where you can go through various informative topics, provide comments, communicate with Tresata experts using Personal Chat options or Emails, etc. \n\nYou will find like minded, Technology Enthusiasts, Data Champions, Tresata Product Experts, and Subject Matter Experts on this Tresata Community. \n\nKnow about using the portal here:\n![image|690x329](upload://n72U8QITc9VRqqzBs68ZRcAgwT5.png)\n\n\n\n\n\n\nYou will see personalised cards displayed on the [landing page](https://community.tresata.com/) covering multiple topic categories with relevant posts, specifically for you. The **GET STARTED** section will help you use the downloaded product easily.\n\nYou can leverage the robust **Search** functionality to find topic you are interested and leave comments, vote for the topic, or even create a new topic if needed.\n\nFor any support required, do reach out to support@tresata.com|false|true|true|4|Welcome to Tresata Community!|4



